`timescale 1ns / 1ps
// Verilog
// c432
// Ninputs 36
// Noutputs 7
// NtotalGates 160
// NOT1 40
// NAND2 64
// NOR2 19
// AND9 3
// XOR2 18
// NAND4 14
// AND8 1
// NAND3 1

module top (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
                  N430,N431,N432,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
                  keyinput30, keyinput31,
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36,
        keyinput37, keyinput38, keyinput39, keyinput40, keyinput41,
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46,
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51,
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56,
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61,
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66,
        keyinput67, keyinput68, keyinput69, keyinput70, keyinput71,
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76,
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81,
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86,
        keyinput87, keyinput88, keyinput89, keyinput90, keyinput91,
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96,
        keyinput97, keyinput98, keyinput99, keyinput100, keyinput101,
                  keyinput102, keyinput103,
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
        keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
        keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
        keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
        keyinput139);

  input keyinput104, keyinput105, keyinput106, keyinput107, keyinput108;
  input keyinput109, keyinput110, keyinput111, keyinput112, keyinput113;
  input keyinput114, keyinput115, keyinput116, keyinput117, keyinput118;
  input keyinput119, keyinput120, keyinput121, keyinput122, keyinput123;
  input keyinput124, keyinput125, keyinput126, keyinput127, keyinput128;
  input keyinput129, keyinput130, keyinput131, keyinput132, keyinput133;
  input keyinput134, keyinput135, keyinput136, keyinput137, keyinput138;
  input keyinput139;


  input keyinput32, keyinput33, keyinput34, keyinput35, keyinput36;
  input keyinput37, keyinput38, keyinput39, keyinput40, keyinput41;
  input keyinput42, keyinput43, keyinput44, keyinput45, keyinput46;
  input keyinput47, keyinput48, keyinput49, keyinput50, keyinput51;
  input keyinput52, keyinput53, keyinput54, keyinput55, keyinput56;
  input keyinput57, keyinput58, keyinput59, keyinput60, keyinput61;
  input keyinput62, keyinput63, keyinput64, keyinput65, keyinput66;
  input keyinput67, keyinput68, keyinput69, keyinput70, keyinput71;
  input keyinput72, keyinput73, keyinput74, keyinput75, keyinput76;
  input keyinput77, keyinput78, keyinput79, keyinput80, keyinput81;
  input keyinput82, keyinput83, keyinput84, keyinput85, keyinput86;
  input keyinput87, keyinput88, keyinput89, keyinput90, keyinput91;
  input keyinput92, keyinput93, keyinput94, keyinput95, keyinput96;
  input keyinput97, keyinput98, keyinput99, keyinput100, keyinput101;
  input keyinput102, keyinput103;

  wire KeyWire_0_1 , KeyWire_0_2;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31;

  wire [0:31] keyinput_Wire_0;
  wire [0:13] KeyNOTWire_0;

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;

output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429;

not NOT1_1 (N118, N1);
not NOT1_2 (N119, N4);
not NOT1_3 (N122, N11);
not NOT1_4 (N123, N17);
  not NOT1_5 (keyinput_Wire_0[0], N24);
  xor keyGate_0_0(KeyNOTWire_0[0], keyinput0, keyinput_Wire_0[0]);
  not KeyNOTGate_0_0(N126, KeyNOTWire_0[0]);
not NOT1_6 (N127, N30);
not NOT1_7 (N130, N37);
not NOT1_8 (N131, N43);
not NOT1_9 (N134, N50);
not NOT1_10 (N135, N56);
not NOT1_11 (N138, N63);
not NOT1_12 (N139, N69);
not NOT1_13 (N142, N76);
not NOT1_14 (N143, N82);
not NOT1_15 (N146, N89);
not NOT1_16 (N147, N95);
  not NOT1_17 (keyinput_Wire_0[1], N102);
  xnor keyGate_0_1(KeyNOTWire_0[1], keyinput1, keyinput_Wire_0[1]);
  not KeyNOTGate_0_1(N150, KeyNOTWire_0[1]);
not NOT1_18 (N151, N108);
nand NAND2_19 (N154, N118, N4);
nor NOR2_20 (N157, N8, N119);
nor NOR2_21 (N158, N14, N119);
nand NAND2_22 (N159, N122, N17);
nand NAND2_23 (N162, N126, N30);
  nand NAND2_24 (keyinput_Wire_0[2], N130, N43);
  xor keyGate_0_2(KeyNOTWire_0[2], keyinput2, keyinput_Wire_0[2]);
  not KeyNOTGate_0_2(N165, KeyNOTWire_0[2]);
  nand NAND2_25 (keyinput_Wire_0[3], N134, N56);
  xor keyGate_0_3(N168, keyinput3, keyinput_Wire_0[3]);
nand NAND2_26 (N171, N138, N69);
nand NAND2_27 (N174, N142, N82);
nand NAND2_28 (N177, N146, N95);
nand NAND2_29 (N180, N150, N108);
nor NOR2_30 (N183, N21, N123);
  nor NOR2_31 (keyinput_Wire_0[4], N27, N123);
  xnor keyGate_0_4(KeyNOTWire_0[3], keyinput4, keyinput_Wire_0[4]);
  not KeyNOTGate_0_3(N184, KeyNOTWire_0[3]);
nor NOR2_32 (N185, N34, N127);
nor NOR2_33 (N186, N40, N127);
nor NOR2_34 (N187, N47, N131);
nor NOR2_35 (N188, N53, N131);
nor NOR2_36 (N189, N60, N135);
nor NOR2_37 (N190, N66, N135);
nor NOR2_38 (N191, N73, N139);
  nor NOR2_39 (keyinput_Wire_0[5], N79, N139);
  xnor keyGate_0_5(N192, keyinput5, keyinput_Wire_0[5]);
nor NOR2_40 (N193, N86, N143);
  nor NOR2_41 (keyinput_Wire_0[6], N92, N143);
  xor keyGate_0_6(KeyNOTWire_0[4], keyinput6, keyinput_Wire_0[6]);
  not KeyNOTGate_0_4(N194, KeyNOTWire_0[4]);
nor NOR2_42 (N195, N99, N147);
nor NOR2_43 (N196, N105, N147);
nor NOR2_44 (N197, N112, N151);
  nor NOR2_45 (keyinput_Wire_0[7], N115, N151);
  xnor keyGate_0_7(N198, keyinput7, keyinput_Wire_0[7]);
  and AND9_46 (keyinput_Wire_0[8], N154, N159, N162, N165, N168, N171, N174, N177, N180);
  xor keyGate_0_8(KeyNOTWire_0[5], keyinput8, keyinput_Wire_0[8]);
  not KeyNOTGate_0_5(N199, KeyNOTWire_0[5]);
not NOT1_47 (N203, N199);
not NOT1_48 (N213, N199);
not NOT1_49 (KeyWire_0_1, N199);
  xor flip_it (N223, KeyWire_0_1, KeyWire_0_2 );
xor XOR2_50 (N224, N203, N154);
xor XOR2_51 (N227, N203, N159);
xor XOR2_52 (N230, N203, N162);
xor XOR2_53 (N233, N203, N165);
xor XOR2_54 (N236, N203, N168);
xor XOR2_55 (N239, N203, N171);
nand NAND2_56 (N242, N1, N213);
xor XOR2_57 (N243, N203, N174);
nand NAND2_58 (N246, N213, N11);
xor XOR2_59 (N247, N203, N177);
  nand NAND2_60 (keyinput_Wire_0[9], N213, N24);
  xnor keyGate_0_9(N250, keyinput9, keyinput_Wire_0[9]);
xor XOR2_61 (N251, N203, N180);
nand NAND2_62 (N254, N213, N37);
nand NAND2_63 (N255, N213, N50);
nand NAND2_64 (N256, N213, N63);
  nand NAND2_65 (keyinput_Wire_0[10], N213, N76);
  xnor keyGate_0_10(N257, keyinput10, keyinput_Wire_0[10]);
  nand NAND2_66 (keyinput_Wire_0[11], N213, N89);
  xnor keyGate_0_11(KeyNOTWire_0[6], keyinput11, keyinput_Wire_0[11]);
  not KeyNOTGate_0_6(N258, KeyNOTWire_0[6]);
  nand NAND2_67 (keyinput_Wire_0[12], N213, N102);
  xor keyGate_0_12(KeyNOTWire_0[7], keyinput12, keyinput_Wire_0[12]);
  not KeyNOTGate_0_7(N259, KeyNOTWire_0[7]);
nand NAND2_68 (N260, N224, N157);
nand NAND2_69 (N263, N224, N158);
nand NAND2_70 (N264, N227, N183);
nand NAND2_71 (N267, N230, N185);
  nand NAND2_72 (keyinput_Wire_0[13], N233, N187);
  xor keyGate_0_13(KeyNOTWire_0[8], keyinput13, keyinput_Wire_0[13]);
  not KeyNOTGate_0_8(N270, KeyNOTWire_0[8]);
  nand NAND2_73 (keyinput_Wire_0[14], N236, N189);
  xnor keyGate_0_14(KeyNOTWire_0[9], keyinput14, keyinput_Wire_0[14]);
  not KeyNOTGate_0_9(N273, KeyNOTWire_0[9]);
nand NAND2_74 (N276, N239, N191);
nand NAND2_75 (N279, N243, N193);
nand NAND2_76 (N282, N247, N195);
nand NAND2_77 (N285, N251, N197);
nand NAND2_78 (N288, N227, N184);
nand NAND2_79 (N289, N230, N186);
nand NAND2_80 (N290, N233, N188);
  nand NAND2_81 (keyinput_Wire_0[15], N236, N190);
  xor keyGate_0_15(KeyNOTWire_0[10], keyinput15, keyinput_Wire_0[15]);
  not KeyNOTGate_0_10(N291, KeyNOTWire_0[10]);
  nand NAND2_82 (keyinput_Wire_0[16], N239, N192);
  xnor keyGate_0_16(N292, keyinput16, keyinput_Wire_0[16]);
nand NAND2_83 (N293, N243, N194);
nand NAND2_84 (N294, N247, N196);
  nand NAND2_85 (keyinput_Wire_0[17], N251, N198);
  xnor keyGate_0_17(N295, keyinput17, keyinput_Wire_0[17]);
and AND9_86 (N296, N260, N264, N267, N270, N273, N276, N279, N282, N285);
not NOT1_87 (N300, N263);
not NOT1_88 (N301, N288);
not NOT1_89 (N302, N289);
not NOT1_90 (N303, N290);
not NOT1_91 (N304, N291);
not NOT1_92 (N305, N292);
not NOT1_93 (N306, N293);
not NOT1_94 (N307, N294);
not NOT1_95 (N308, N295);
  not NOT1_96 (keyinput_Wire_0[18], N296);
  xor keyGate_0_18(N309, keyinput18, keyinput_Wire_0[18]);
not NOT1_97 (N319, N296);
not NOT1_98 (N329, N296);
xor XOR2_99 (N330, N309, N260);
xor XOR2_100 (N331, N309, N264);
xor XOR2_101 (N332, N309, N267);
xor XOR2_102 (N333, N309, N270);
nand NAND2_103 (N334, N8, N319);
xor XOR2_104 (N335, N309, N273);
nand NAND2_105 (N336, N319, N21);
xor XOR2_106 (N337, N309, N276);
nand NAND2_107 (N338, N319, N34);
  xor XOR2_108 (keyinput_Wire_0[19], N309, N279);
  xor keyGate_0_19(N339, keyinput19, keyinput_Wire_0[19]);
  nand NAND2_109 (keyinput_Wire_0[20], N319, N47);
  xor keyGate_0_20(KeyNOTWire_0[11], keyinput20, keyinput_Wire_0[20]);
  not KeyNOTGate_0_11(N340, KeyNOTWire_0[11]);
xor XOR2_110 (N341, N309, N282);
nand NAND2_111 (N342, N319, N60);
xor XOR2_112 (N343, N309, N285);
nand NAND2_113 (N344, N319, N73);
nand NAND2_114 (N345, N319, N86);
nand NAND2_115 (N346, N319, N99);
nand NAND2_116 (N347, N319, N112);
nand NAND2_117 (N348, N330, N300);
nand NAND2_118 (N349, N331, N301);
nand NAND2_119 (N350, N332, N302);
  nand NAND2_120 (keyinput_Wire_0[21], N333, N303);
  xnor keyGate_0_21(N351, keyinput21, keyinput_Wire_0[21]);
nand NAND2_121 (N352, N335, N304);
nand NAND2_122 (N353, N337, N305);
nand NAND2_123 (N354, N339, N306);
nand NAND2_124 (N355, N341, N307);
nand NAND2_125 (N356, N343, N308);
and AND9_126 (N357, N348, N349, N350, N351, N352, N353, N354, N355, N356);
not NOT1_127 (N360, N357);
not NOT1_128 (N370, N357);
nand NAND2_129 (N371, N14, N360);
  nand NAND2_130 (keyinput_Wire_0[22], N360, N27);
  xnor keyGate_0_22(KeyNOTWire_0[12], keyinput22, keyinput_Wire_0[22]);
  not KeyNOTGate_0_12(N372, KeyNOTWire_0[12]);
nand NAND2_131 (N373, N360, N40);
nand NAND2_132 (N374, N360, N53);
nand NAND2_133 (N375, N360, N66);
  nand NAND2_134 (keyinput_Wire_0[23], N360, N79);
  xnor keyGate_0_23(N376, keyinput23, keyinput_Wire_0[23]);
  nand NAND2_135 (keyinput_Wire_0[24], N360, N92);
  xnor keyGate_0_24(N377, keyinput24, keyinput_Wire_0[24]);
nand NAND2_136 (N378, N360, N105);
nand NAND2_137 (N379, N360, N115);
nand NAND4_138 (N380, N4, N242, N334, N371);
nand NAND4_139 (N381, N246, N336, N372, N17);
nand NAND4_140 (N386, N250, N338, N373, N30);
  nand NAND4_141 (keyinput_Wire_0[25], N254, N340, N374, N43);
  xor keyGate_0_25(N393, keyinput25, keyinput_Wire_0[25]);
nand NAND4_142 (N399, N255, N342, N375, N56);
nand NAND4_143 (N404, N256, N344, N376, N69);
nand NAND4_144 (N407, N257, N345, N377, N82);
nand NAND4_145 (N411, N258, N346, N378, N95);
  nand NAND4_146 (keyinput_Wire_0[26], N259, N347, N379, N108);
  xor keyGate_0_26(N414, keyinput26, keyinput_Wire_0[26]);
  not NOT1_147 (keyinput_Wire_0[27], N380);
  xnor keyGate_0_27(KeyNOTWire_0[13], keyinput27, keyinput_Wire_0[27]);
  not KeyNOTGate_0_13(N415, KeyNOTWire_0[13]);
  and AND8_148 (keyinput_Wire_0[28], N381, N386, N393, N399, N404, N407, N411, N414);
  xnor keyGate_0_28(N416, keyinput28, keyinput_Wire_0[28]);
not NOT1_149 (N417, N393);
not NOT1_150 (N418, N404);
not NOT1_151 (N419, N407);
  not NOT1_152 (keyinput_Wire_0[29], N411);
  xor keyGate_0_29(N420, keyinput29, keyinput_Wire_0[29]);
nor NOR2_153 (N421, N415, N416);
  nand NAND2_154 (keyinput_Wire_0[30], N386, N417);
  xor keyGate_0_30(N422, keyinput30, keyinput_Wire_0[30]);
nand NAND4_155 (N425, N386, N393, N418, N399);
  nand NAND3_156 (keyinput_Wire_0[31], N399, N393, N419);
  xnor keyGate_0_31(N428, keyinput31, keyinput_Wire_0[31]);
nand NAND4_157 (N429, N386, N393, N407, N420);
nand NAND4_158 (N430, N381, N386, N422, N399);
nand NAND4_159 (N431, N381, N386, N425, N428);
nand NAND4_160 (N432, N381, N422, N425, N429);

AntiSAT some_name( KeyWire_0_2, N115, N63, N43, N1, N8, N47, N27, N14, N53, N17, N69, N11, N60, N112, N40, N50, N108, N82, N66, N21, N30, N105, N76, N73, N4, N102, N89, N24, N99, N79, N34, N95, N56, N37, N86, N92, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
       keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
       keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
       keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
       keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
       keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
       keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
       keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
       keyinput139);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N115, N63, N43, N1, N8, N47, N27, N14, N53, N17, N69, N11, N60, N112, N40, N50, N108, N82, N66, N21, N30, N105, N76, N73, N4, N102, N89, N24, N99, N79, N34, N95, N56, N37, N86, N92, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103 ,
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
        keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
        keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
        keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
        keyinput139);

  input keyinput104, keyinput105, keyinput106, keyinput107, keyinput108;
  input keyinput109, keyinput110, keyinput111, keyinput112, keyinput113;
  input keyinput114, keyinput115, keyinput116, keyinput117, keyinput118;
  input keyinput119, keyinput120, keyinput121, keyinput122, keyinput123;
  input keyinput124, keyinput125, keyinput126, keyinput127, keyinput128;
  input keyinput129, keyinput130, keyinput131, keyinput132, keyinput133;
  input keyinput134, keyinput135, keyinput136, keyinput137, keyinput138;
  input keyinput139;

  wire [0:35] keyNTin_Wire_1;
  wire [0:13] KeyNOTWire_1;

  input N115, N63, N43, N1, N8, N47, N27, N14, N53, N17, N69, N11, N60, N112, N40, N50, N108, N82, N66, N21, N30, N105, N76, N73, N4, N102, N89, N24, N99, N79, N34, N95, N56, N37, N86, N92;
  input keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73 ;

  xnor KeyGate0 (keyNTin_Wire_1[0], N115, keyinput32);
  xor keyNTinGate_1_0(newWire_0, keyinput104, keyNTin_Wire_1[0]);
  xnor KeyGate1 (keyNTin_Wire_1[1], N63, keyinput33);
  xor keyNTinGate_1_1(newWire_1, keyinput105, keyNTin_Wire_1[1]);
  xnor KeyGate2 (keyNTin_Wire_1[2], N43, keyinput34);
  xor keyNTinGate_1_2(newWire_2, keyinput106, keyNTin_Wire_1[2]);
  xor  KeyGate3 (newWire_3, N1, keyinput35);
  xnor KeyGate4 (keyNTin_Wire_1[3], N8, keyinput36);
  xnor keyNTinGate_1_3(newWire_4, keyinput107, keyNTin_Wire_1[3]);
  xor  KeyGate5 (keyNTin_Wire_1[4], N47, keyinput37);
  xor keyNTinGate_1_4(newWire_5, keyinput108, keyNTin_Wire_1[4]);
  xor  KeyGate6 (keyNTin_Wire_1[5], N27, keyinput38);
  xnor keyNTinGate_1_5(KeyNOTWire_1[0], keyinput109, keyNTin_Wire_1[5]);
  not KeyNOTGate_1_0(newWire_6, KeyNOTWire_1[0]);
  xor  KeyGate7 (keyNTin_Wire_1[6], N14, keyinput39);
  xnor keyNTinGate_1_6(newWire_7, keyinput110, keyNTin_Wire_1[6]);
  xor  KeyGate8 (keyNTin_Wire_1[7], N53, keyinput40);
  xnor keyNTinGate_1_7(newWire_8, keyinput111, keyNTin_Wire_1[7]);
  xor  KeyGate9 (keyNTin_Wire_1[8], N17, keyinput41);
  xnor keyNTinGate_1_8(KeyNOTWire_1[1], keyinput112, keyNTin_Wire_1[8]);
  not KeyNOTGate_1_1(newWire_9, KeyNOTWire_1[1]);
  xnor KeyGate10 (keyNTin_Wire_1[9], N69, keyinput42);
  xor keyNTinGate_1_9(newWire_10, keyinput113, keyNTin_Wire_1[9]);
  xnor KeyGate11 (keyNTin_Wire_1[10], N11, keyinput43);
  xnor keyNTinGate_1_10(KeyNOTWire_1[2], keyinput114, keyNTin_Wire_1[10]);
  not KeyNOTGate_1_2(newWire_11, KeyNOTWire_1[2]);
  xnor KeyGate12 (keyNTin_Wire_1[11], N60, keyinput44);
  xor keyNTinGate_1_11(newWire_12, keyinput115, keyNTin_Wire_1[11]);
  xor  KeyGate13 (keyNTin_Wire_1[12], N112, keyinput45);
  xor keyNTinGate_1_12(KeyNOTWire_1[3], keyinput116, keyNTin_Wire_1[12]);
  not KeyNOTGate_1_3(newWire_13, KeyNOTWire_1[3]);
  xor  KeyGate14 (newWire_14, N40, keyinput46);
  xor  KeyGate15 (keyNTin_Wire_1[13], N50, keyinput47);
  xor keyNTinGate_1_13(KeyNOTWire_1[4], keyinput117, keyNTin_Wire_1[13]);
  not KeyNOTGate_1_4(newWire_15, KeyNOTWire_1[4]);
  xnor KeyGate16 (keyNTin_Wire_1[14], N108, keyinput48);
  xnor keyNTinGate_1_14(newWire_16, keyinput118, keyNTin_Wire_1[14]);
  xor  KeyGate17 (keyNTin_Wire_1[15], N82, keyinput49);
  xnor keyNTinGate_1_15(KeyNOTWire_1[5], keyinput119, keyNTin_Wire_1[15]);
  not KeyNOTGate_1_5(newWire_17, KeyNOTWire_1[5]);
  xnor KeyGate18 (keyNTin_Wire_1[16], N66, keyinput50);
  xnor keyNTinGate_1_16(newWire_18, keyinput120, keyNTin_Wire_1[16]);
  xnor KeyGate19 (newWire_19, N21, keyinput51);
  xnor KeyGate20 (newWire_20, N30, keyinput52);
  xor  KeyGate21 (newWire_21, N105, keyinput53);
  xnor KeyGate22 (keyNTin_Wire_1[17], N76, keyinput54);
  xnor keyNTinGate_1_17(newWire_22, keyinput121, keyNTin_Wire_1[17]);
  xor  KeyGate23 (newWire_23, N73, keyinput55);
  xnor KeyGate24 (newWire_24, N4, keyinput56);
  xor  KeyGate25 (keyNTin_Wire_1[18], N102, keyinput57);
  xor keyNTinGate_1_18(newWire_25, keyinput122, keyNTin_Wire_1[18]);
  xnor KeyGate26 (newWire_26, N89, keyinput58);
  xnor KeyGate27 (keyNTin_Wire_1[19], N24, keyinput59);
  xor keyNTinGate_1_19(newWire_27, keyinput123, keyNTin_Wire_1[19]);
  xor  KeyGate28 (newWire_28, N99, keyinput60);
  xnor KeyGate29 (newWire_29, N79, keyinput61);
  xor  KeyGate30 (newWire_30, N34, keyinput62);
  xor  KeyGate31 (newWire_31, N95, keyinput63);
  xor  KeyGate32 (newWire_32, N56, keyinput64);
  xor  KeyGate33 (newWire_33, N37, keyinput65);
  xnor KeyGate34 (keyNTin_Wire_1[20], N86, keyinput66);
  xnor keyNTinGate_1_20(KeyNOTWire_1[6], keyinput124, keyNTin_Wire_1[20]);
  not KeyNOTGate_1_6(newWire_34, KeyNOTWire_1[6]);
  xor  KeyGate35 (newWire_35, N92, keyinput67);
  xnor KeyGate36 (keyNTin_Wire_1[21], N115, keyinput68);
  xnor keyNTinGate_1_21(newWire_36, keyinput125, keyNTin_Wire_1[21]);
  xnor KeyGate37 (newWire_37, N63, keyinput69);
  xor  KeyGate38 (keyNTin_Wire_1[22], N43, keyinput70);
  xor keyNTinGate_1_22(KeyNOTWire_1[7], keyinput126, keyNTin_Wire_1[22]);
  not KeyNOTGate_1_7(newWire_38, KeyNOTWire_1[7]);
  xnor KeyGate39 (newWire_39, N1, keyinput71);
  xnor KeyGate40 (newWire_40, N8, keyinput72);
  xor  KeyGate41 (newWire_41, N47, keyinput73);
  xor  KeyGate42 (newWire_42, N27, keyinput74);
  xnor KeyGate43 (newWire_43, N14, keyinput75);
  xor  KeyGate44 (newWire_44, N53, keyinput76);
  xor  KeyGate45 (keyNTin_Wire_1[23], N17, keyinput77);
  xor keyNTinGate_1_23(KeyNOTWire_1[8], keyinput127, keyNTin_Wire_1[23]);
  not KeyNOTGate_1_8(newWire_45, KeyNOTWire_1[8]);
  xor  KeyGate46 (keyNTin_Wire_1[24], N69, keyinput78);
  xnor keyNTinGate_1_24(KeyNOTWire_1[9], keyinput128, keyNTin_Wire_1[24]);
  not KeyNOTGate_1_9(newWire_46, KeyNOTWire_1[9]);
  xnor KeyGate47 (newWire_47, N11, keyinput79);
  xor  KeyGate48 (newWire_48, N60, keyinput80);
  xor  KeyGate49 (newWire_49, N112, keyinput81);
  xor  KeyGate50 (newWire_50, N40, keyinput82);
  xnor KeyGate51 (newWire_51, N50, keyinput83);
  xor  KeyGate52 (keyNTin_Wire_1[25], N108, keyinput84);
  xnor keyNTinGate_1_25(newWire_52, keyinput129, keyNTin_Wire_1[25]);
  xnor KeyGate53 (newWire_53, N82, keyinput85);
  xnor KeyGate54 (newWire_54, N66, keyinput86);
  xnor KeyGate55 (newWire_55, N21, keyinput87);
  xnor KeyGate56 (newWire_56, N30, keyinput88);
  xnor KeyGate57 (newWire_57, N105, keyinput89);
  xnor KeyGate58 (keyNTin_Wire_1[26], N76, keyinput90);
  xnor keyNTinGate_1_26(KeyNOTWire_1[10], keyinput130, keyNTin_Wire_1[26]);
  not KeyNOTGate_1_10(newWire_58, KeyNOTWire_1[10]);
  xor  KeyGate59 (newWire_59, N73, keyinput91);
  xor  KeyGate60 (keyNTin_Wire_1[27], N4, keyinput92);
  xor keyNTinGate_1_27(KeyNOTWire_1[11], keyinput131, keyNTin_Wire_1[27]);
  not KeyNOTGate_1_11(newWire_60, KeyNOTWire_1[11]);
  xnor KeyGate61 (newWire_61, N102, keyinput93);
  xnor KeyGate62 (keyNTin_Wire_1[28], N89, keyinput94);
  xnor keyNTinGate_1_28(newWire_62, keyinput132, keyNTin_Wire_1[28]);
  xnor KeyGate63 (newWire_63, N24, keyinput95);
  xnor KeyGate64 (newWire_64, N99, keyinput96);
  xor  KeyGate65 (newWire_65, N79, keyinput97);
  xnor KeyGate66 (keyNTin_Wire_1[29], N34, keyinput98);
  xor keyNTinGate_1_29(newWire_66, keyinput133, keyNTin_Wire_1[29]);
  xor  KeyGate67 (keyNTin_Wire_1[30], N95, keyinput99);
  xor keyNTinGate_1_30(newWire_67, keyinput134, keyNTin_Wire_1[30]);
  xnor KeyGate68 (keyNTin_Wire_1[31], N56, keyinput100);
  xnor keyNTinGate_1_31(newWire_68, keyinput135, keyNTin_Wire_1[31]);
  xnor KeyGate69 (keyNTin_Wire_1[32], N37, keyinput101);
  xor keyNTinGate_1_32(KeyNOTWire_1[12], keyinput136, keyNTin_Wire_1[32]);
  not KeyNOTGate_1_12(newWire_69, KeyNOTWire_1[12]);
  xnor KeyGate70 (newWire_70, N86, keyinput102);
  xnor KeyGate71 (keyNTin_Wire_1[33], N92, keyinput103);
  xnor keyNTinGate_1_33(newWire_71, keyinput137, keyNTin_Wire_1[33]);
  and some_function (newWire_72, newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35 );
  nand compl_function (keyNTin_Wire_1[34], newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71);
  xnor keyNTinGate_1_34(KeyNOTWire_1[13], keyinput138, keyNTin_Wire_1[34]);
  not KeyNOTGate_1_13(newWire_73, KeyNOTWire_1[13]);
  and finalAND (keyNTin_Wire_1[35], newWire_72, newWire_73);
  xor keyNTinGate_1_35(KeyWire_0_2, keyinput139, keyNTin_Wire_1[35]);

endmodule /* AntiSAT */
