`timescale 1ns / 1ps
// Verilog
// c880
// Ninputs 60
// Noutputs 26
// NtotalGates 383
// NAND4 13
// AND3 12
// NAND2 60
// NAND3 14
// AND2 105
// OR2 29
// NOT1 63
// NOR2 61
// BUFF1 26

module top (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
                  N865,N866,N874,N878,N879,N880,
        keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4,
        keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9,
        keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14,
        keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19,
        keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24,
        keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29,
        keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34,
        keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39,
        keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44,
        keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49,
        keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54,
        keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59,
        keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64,
        keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69,
        keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74,
        keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79,
        keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84,
        keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89,
        keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94,
        keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99,
        keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104,
        keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109,
        keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114,
        keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119,
        keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124,
        keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129,
        keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134,
        keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139,
        keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144,
        keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149,
        keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154,
        keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159,
        keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164,
        keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169,
        keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174,
        keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179,
        keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184,
        keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189,
        keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194,
        keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199,
        keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204,
        keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209,
        keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214,
        keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219,
        keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224,
        keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229,
        keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234,
        keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239,
        keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244,
        keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249,
        keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254,
        keyIn_0_255);

  input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4;
  input keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9;
  input keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14;
  input keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19;
  input keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24;
  input keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29;
  input keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34;
  input keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39;
  input keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44;
  input keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49;
  input keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54;
  input keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59;
  input keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64;
  input keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69;
  input keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74;
  input keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79;
  input keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84;
  input keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89;
  input keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94;
  input keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99;
  input keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104;
  input keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109;
  input keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114;
  input keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119;
  input keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124;
  input keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129;
  input keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134;
  input keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139;
  input keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144;
  input keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149;
  input keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154;
  input keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159;
  input keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164;
  input keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169;
  input keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174;
  input keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179;
  input keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184;
  input keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189;
  input keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194;
  input keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199;
  input keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204;
  input keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209;
  input keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214;
  input keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219;
  input keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224;
  input keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229;
  input keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234;
  input keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239;
  input keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244;
  input keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249;
  input keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254;
  input keyIn_0_255;

  wire [0:255] KeyWire_0;
  wire [0:125] KeyNOTWire_0;

input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;

output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;

wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877;

  nand NAND4_1 (KeyWire_0[0], N1, N8, N13, N17);
  xnor KeyGate_0_0(KeyNOTWire_0[0], keyIn_0_0, KeyWire_0[0]);
  not KeyNOTGate_0_0(N269, KeyNOTWire_0[0]);
  nand NAND4_2 (KeyWire_0[1], N1, N26, N13, N17);
  xnor KeyGate_0_1(N270, keyIn_0_1, KeyWire_0[1]);
  and AND3_3 (KeyWire_0[2], N29, N36, N42);
  xor KeyGate_0_2(N273, keyIn_0_2, KeyWire_0[2]);
and AND3_4 (N276, N1, N26, N51);
  nand NAND4_5 (KeyWire_0[3], N1, N8, N51, N17);
  xor KeyGate_0_3(N279, keyIn_0_3, KeyWire_0[3]);
nand NAND4_6 (N280, N1, N8, N13, N55);
  nand NAND4_7 (KeyWire_0[4], N59, N42, N68, N72);
  xnor KeyGate_0_4(KeyNOTWire_0[1], keyIn_0_4, KeyWire_0[4]);
  not KeyNOTGate_0_1(N284, KeyNOTWire_0[1]);
nand NAND2_8 (N285, N29, N68);
nand NAND3_9 (N286, N59, N68, N74);
and AND3_10 (N287, N29, N75, N80);
  and AND3_11 (KeyWire_0[5], N29, N75, N42);
  xnor KeyGate_0_5(KeyNOTWire_0[2], keyIn_0_5, KeyWire_0[5]);
  not KeyNOTGate_0_2(N290, KeyNOTWire_0[2]);
  and AND3_12 (KeyWire_0[6], N29, N36, N80);
  xor KeyGate_0_6(N291, keyIn_0_6, KeyWire_0[6]);
and AND3_13 (N292, N29, N36, N42);
  and AND3_14 (KeyWire_0[7], N59, N75, N80);
  xor KeyGate_0_7(N293, keyIn_0_7, KeyWire_0[7]);
  and AND3_15 (KeyWire_0[8], N59, N75, N42);
  xor KeyGate_0_8(KeyNOTWire_0[3], keyIn_0_8, KeyWire_0[8]);
  not KeyNOTGate_0_3(N294, KeyNOTWire_0[3]);
  and AND3_16 (KeyWire_0[9], N59, N36, N80);
  xnor KeyGate_0_9(N295, keyIn_0_9, KeyWire_0[9]);
  and AND3_17 (KeyWire_0[10], N59, N36, N42);
  xnor KeyGate_0_10(N296, keyIn_0_10, KeyWire_0[10]);
  and AND2_18 (KeyWire_0[11], N85, N86);
  xnor KeyGate_0_11(KeyNOTWire_0[4], keyIn_0_11, KeyWire_0[11]);
  not KeyNOTGate_0_4(N297, KeyNOTWire_0[4]);
  or OR2_19 (KeyWire_0[12], N87, N88);
  xnor KeyGate_0_12(N298, keyIn_0_12, KeyWire_0[12]);
  nand NAND2_20 (KeyWire_0[13], N91, N96);
  xnor KeyGate_0_13(N301, keyIn_0_13, KeyWire_0[13]);
  or OR2_21 (KeyWire_0[14], N91, N96);
  xor KeyGate_0_14(N302, keyIn_0_14, KeyWire_0[14]);
nand NAND2_22 (N303, N101, N106);
  or OR2_23 (KeyWire_0[15], N101, N106);
  xor KeyGate_0_15(N304, keyIn_0_15, KeyWire_0[15]);
  nand NAND2_24 (KeyWire_0[16], N111, N116);
  xor KeyGate_0_16(N305, keyIn_0_16, KeyWire_0[16]);
  or OR2_25 (KeyWire_0[17], N111, N116);
  xor KeyGate_0_17(KeyNOTWire_0[5], keyIn_0_17, KeyWire_0[17]);
  not KeyNOTGate_0_5(N306, KeyNOTWire_0[5]);
nand NAND2_26 (N307, N121, N126);
  or OR2_27 (KeyWire_0[18], N121, N126);
  xnor KeyGate_0_18(KeyNOTWire_0[6], keyIn_0_18, KeyWire_0[18]);
  not KeyNOTGate_0_6(N308, KeyNOTWire_0[6]);
and AND2_28 (N309, N8, N138);
  not NOT1_29 (KeyWire_0[19], N268);
  xnor KeyGate_0_19(KeyNOTWire_0[7], keyIn_0_19, KeyWire_0[19]);
  not KeyNOTGate_0_7(N310, KeyNOTWire_0[7]);
  and AND2_30 (KeyWire_0[20], N51, N138);
  xnor KeyGate_0_20(N316, keyIn_0_20, KeyWire_0[20]);
  and AND2_31 (KeyWire_0[21], N17, N138);
  xnor KeyGate_0_21(KeyNOTWire_0[8], keyIn_0_21, KeyWire_0[21]);
  not KeyNOTGate_0_8(N317, KeyNOTWire_0[8]);
and AND2_32 (N318, N152, N138);
  nand NAND2_33 (KeyWire_0[22], N59, N156);
  xor KeyGate_0_22(N319, keyIn_0_22, KeyWire_0[22]);
  nor NOR2_34 (KeyWire_0[23], N17, N42);
  xor KeyGate_0_23(KeyNOTWire_0[9], keyIn_0_23, KeyWire_0[23]);
  not KeyNOTGate_0_9(N322, KeyNOTWire_0[9]);
  and AND2_35 (KeyWire_0[24], N17, N42);
  xor KeyGate_0_24(N323, keyIn_0_24, KeyWire_0[24]);
  nand NAND2_36 (KeyWire_0[25], N159, N165);
  xor KeyGate_0_25(KeyNOTWire_0[10], keyIn_0_25, KeyWire_0[25]);
  not KeyNOTGate_0_10(N324, KeyNOTWire_0[10]);
  or OR2_37 (KeyWire_0[26], N159, N165);
  xor KeyGate_0_26(N325, keyIn_0_26, KeyWire_0[26]);
  nand NAND2_38 (KeyWire_0[27], N171, N177);
  xnor KeyGate_0_27(KeyNOTWire_0[11], keyIn_0_27, KeyWire_0[27]);
  not KeyNOTGate_0_11(N326, KeyNOTWire_0[11]);
  or OR2_39 (KeyWire_0[28], N171, N177);
  xor KeyGate_0_28(KeyNOTWire_0[12], keyIn_0_28, KeyWire_0[28]);
  not KeyNOTGate_0_12(N327, KeyNOTWire_0[12]);
nand NAND2_40 (N328, N183, N189);
  or OR2_41 (KeyWire_0[29], N183, N189);
  xor KeyGate_0_29(N329, keyIn_0_29, KeyWire_0[29]);
  nand NAND2_42 (KeyWire_0[30], N195, N201);
  xnor KeyGate_0_30(N330, keyIn_0_30, KeyWire_0[30]);
  or OR2_43 (KeyWire_0[31], N195, N201);
  xor KeyGate_0_31(N331, keyIn_0_31, KeyWire_0[31]);
  and AND2_44 (KeyWire_0[32], N210, N91);
  xnor KeyGate_0_32(KeyNOTWire_0[13], keyIn_0_32, KeyWire_0[32]);
  not KeyNOTGate_0_13(N332, KeyNOTWire_0[13]);
  and AND2_45 (KeyWire_0[33], N210, N96);
  xnor KeyGate_0_33(KeyNOTWire_0[14], keyIn_0_33, KeyWire_0[33]);
  not KeyNOTGate_0_14(N333, KeyNOTWire_0[14]);
and AND2_46 (N334, N210, N101);
  and AND2_47 (KeyWire_0[34], N210, N106);
  xor KeyGate_0_34(N335, keyIn_0_34, KeyWire_0[34]);
  and AND2_48 (KeyWire_0[35], N210, N111);
  xnor KeyGate_0_35(KeyNOTWire_0[15], keyIn_0_35, KeyWire_0[35]);
  not KeyNOTGate_0_15(N336, KeyNOTWire_0[15]);
  and AND2_49 (KeyWire_0[36], N255, N259);
  xor KeyGate_0_36(KeyNOTWire_0[16], keyIn_0_36, KeyWire_0[36]);
  not KeyNOTGate_0_16(N337, KeyNOTWire_0[16]);
and AND2_50 (N338, N210, N116);
  and AND2_51 (KeyWire_0[37], N255, N260);
  xnor KeyGate_0_37(KeyNOTWire_0[17], keyIn_0_37, KeyWire_0[37]);
  not KeyNOTGate_0_17(N339, KeyNOTWire_0[17]);
  and AND2_52 (KeyWire_0[38], N210, N121);
  xnor KeyGate_0_38(KeyNOTWire_0[18], keyIn_0_38, KeyWire_0[38]);
  not KeyNOTGate_0_18(N340, KeyNOTWire_0[18]);
  and AND2_53 (KeyWire_0[39], N255, N267);
  xor KeyGate_0_39(N341, keyIn_0_39, KeyWire_0[39]);
  not NOT1_54 (KeyWire_0[40], N269);
  xor KeyGate_0_40(N342, keyIn_0_40, KeyWire_0[40]);
  not NOT1_55 (KeyWire_0[41], N273);
  xnor KeyGate_0_41(KeyNOTWire_0[19], keyIn_0_41, KeyWire_0[41]);
  not KeyNOTGate_0_19(N343, KeyNOTWire_0[19]);
or OR2_56 (N344, N270, N273);
  not NOT1_57 (KeyWire_0[42], N276);
  xnor KeyGate_0_42(KeyNOTWire_0[20], keyIn_0_42, KeyWire_0[42]);
  not KeyNOTGate_0_20(N345, KeyNOTWire_0[20]);
  not NOT1_58 (KeyWire_0[43], N276);
  xor KeyGate_0_43(KeyNOTWire_0[21], keyIn_0_43, KeyWire_0[43]);
  not KeyNOTGate_0_21(N346, KeyNOTWire_0[21]);
not NOT1_59 (N347, N279);
  nor NOR2_60 (KeyWire_0[44], N280, N284);
  xor KeyGate_0_44(N348, keyIn_0_44, KeyWire_0[44]);
or OR2_61 (N349, N280, N285);
  or OR2_62 (KeyWire_0[45], N280, N286);
  xnor KeyGate_0_45(N350, keyIn_0_45, KeyWire_0[45]);
  not NOT1_63 (KeyWire_0[46], N293);
  xnor KeyGate_0_46(KeyNOTWire_0[22], keyIn_0_46, KeyWire_0[46]);
  not KeyNOTGate_0_22(N351, KeyNOTWire_0[22]);
not NOT1_64 (N352, N294);
  not NOT1_65 (KeyWire_0[47], N295);
  xor KeyGate_0_47(N353, keyIn_0_47, KeyWire_0[47]);
  not NOT1_66 (KeyWire_0[48], N296);
  xor KeyGate_0_48(N354, keyIn_0_48, KeyWire_0[48]);
  nand NAND2_67 (KeyWire_0[49], N89, N298);
  xnor KeyGate_0_49(N355, keyIn_0_49, KeyWire_0[49]);
  and AND2_68 (KeyWire_0[50], N90, N298);
  xnor KeyGate_0_50(KeyNOTWire_0[23], keyIn_0_50, KeyWire_0[50]);
  not KeyNOTGate_0_23(N356, KeyNOTWire_0[23]);
  nand NAND2_69 (KeyWire_0[51], N301, N302);
  xor KeyGate_0_51(N357, keyIn_0_51, KeyWire_0[51]);
nand NAND2_70 (N360, N303, N304);
  nand NAND2_71 (KeyWire_0[52], N305, N306);
  xor KeyGate_0_52(KeyNOTWire_0[24], keyIn_0_52, KeyWire_0[52]);
  not KeyNOTGate_0_24(N363, KeyNOTWire_0[24]);
  nand NAND2_72 (KeyWire_0[53], N307, N308);
  xnor KeyGate_0_53(N366, keyIn_0_53, KeyWire_0[53]);
  not NOT1_73 (KeyWire_0[54], N310);
  xnor KeyGate_0_54(N369, keyIn_0_54, KeyWire_0[54]);
  nor NOR2_74 (KeyWire_0[55], N322, N323);
  xor KeyGate_0_55(KeyNOTWire_0[25], keyIn_0_55, KeyWire_0[55]);
  not KeyNOTGate_0_25(N375, KeyNOTWire_0[25]);
nand NAND2_75 (N376, N324, N325);
nand NAND2_76 (N379, N326, N327);
  nand NAND2_77 (KeyWire_0[56], N328, N329);
  xnor KeyGate_0_56(KeyNOTWire_0[26], keyIn_0_56, KeyWire_0[56]);
  not KeyNOTGate_0_26(N382, KeyNOTWire_0[26]);
  nand NAND2_78 (KeyWire_0[57], N330, N331);
  xor KeyGate_0_57(KeyNOTWire_0[27], keyIn_0_57, KeyWire_0[57]);
  not KeyNOTGate_0_27(N385, KeyNOTWire_0[27]);
buf BUFF1_79 (N388, N290);
buf BUFF1_80 (N389, N291);
buf BUFF1_81 (N390, N292);
buf BUFF1_82 (N391, N297);
  or OR2_83 (KeyWire_0[58], N270, N343);
  xor KeyGate_0_58(N392, keyIn_0_58, KeyWire_0[58]);
  not NOT1_84 (KeyWire_0[59], N345);
  xnor KeyGate_0_59(N393, keyIn_0_59, KeyWire_0[59]);
  not NOT1_85 (KeyWire_0[60], N346);
  xnor KeyGate_0_60(KeyNOTWire_0[28], keyIn_0_60, KeyWire_0[60]);
  not KeyNOTGate_0_28(N399, KeyNOTWire_0[28]);
  and AND2_86 (KeyWire_0[61], N348, N73);
  xor KeyGate_0_61(KeyNOTWire_0[29], keyIn_0_61, KeyWire_0[61]);
  not KeyNOTGate_0_29(N400, KeyNOTWire_0[29]);
  not NOT1_87 (KeyWire_0[62], N349);
  xor KeyGate_0_62(N401, keyIn_0_62, KeyWire_0[62]);
  not NOT1_88 (KeyWire_0[63], N350);
  xnor KeyGate_0_63(KeyNOTWire_0[30], keyIn_0_63, KeyWire_0[63]);
  not KeyNOTGate_0_30(N402, KeyNOTWire_0[30]);
not NOT1_89 (N403, N355);
  not NOT1_90 (KeyWire_0[64], N357);
  xnor KeyGate_0_64(N404, keyIn_0_64, KeyWire_0[64]);
  not NOT1_91 (KeyWire_0[65], N360);
  xor KeyGate_0_65(KeyNOTWire_0[31], keyIn_0_65, KeyWire_0[65]);
  not KeyNOTGate_0_31(N405, KeyNOTWire_0[31]);
  and AND2_92 (KeyWire_0[66], N357, N360);
  xor KeyGate_0_66(N406, keyIn_0_66, KeyWire_0[66]);
  not NOT1_93 (KeyWire_0[67], N363);
  xnor KeyGate_0_67(N407, keyIn_0_67, KeyWire_0[67]);
  not NOT1_94 (KeyWire_0[68], N366);
  xor KeyGate_0_68(KeyNOTWire_0[32], keyIn_0_68, KeyWire_0[68]);
  not KeyNOTGate_0_32(N408, KeyNOTWire_0[32]);
  and AND2_95 (KeyWire_0[69], N363, N366);
  xnor KeyGate_0_69(N409, keyIn_0_69, KeyWire_0[69]);
  nand NAND2_96 (KeyWire_0[70], N347, N352);
  xor KeyGate_0_70(N410, keyIn_0_70, KeyWire_0[70]);
  not NOT1_97 (KeyWire_0[71], N376);
  xor KeyGate_0_71(KeyNOTWire_0[33], keyIn_0_71, KeyWire_0[71]);
  not KeyNOTGate_0_33(N411, KeyNOTWire_0[33]);
  not NOT1_98 (KeyWire_0[72], N379);
  xnor KeyGate_0_72(N412, keyIn_0_72, KeyWire_0[72]);
and AND2_99 (N413, N376, N379);
not NOT1_100 (N414, N382);
  not NOT1_101 (KeyWire_0[73], N385);
  xor KeyGate_0_73(N415, keyIn_0_73, KeyWire_0[73]);
  and AND2_102 (KeyWire_0[74], N382, N385);
  xor KeyGate_0_74(KeyNOTWire_0[34], keyIn_0_74, KeyWire_0[74]);
  not KeyNOTGate_0_34(N416, KeyNOTWire_0[34]);
  and AND2_103 (KeyWire_0[75], N210, N369);
  xnor KeyGate_0_75(N417, keyIn_0_75, KeyWire_0[75]);
buf BUFF1_104 (N418, N342);
buf BUFF1_105 (N419, N344);
buf BUFF1_106 (N420, N351);
buf BUFF1_107 (N421, N353);
buf BUFF1_108 (N422, N354);
buf BUFF1_109 (N423, N356);
  not NOT1_110 (KeyWire_0[76], N400);
  xor KeyGate_0_76(KeyNOTWire_0[35], keyIn_0_76, KeyWire_0[76]);
  not KeyNOTGate_0_35(N424, KeyNOTWire_0[35]);
  and AND2_111 (KeyWire_0[77], N404, N405);
  xor KeyGate_0_77(N425, keyIn_0_77, KeyWire_0[77]);
  and AND2_112 (KeyWire_0[78], N407, N408);
  xor KeyGate_0_78(N426, keyIn_0_78, KeyWire_0[78]);
  and AND3_113 (KeyWire_0[79], N319, N393, N55);
  xor KeyGate_0_79(KeyNOTWire_0[36], keyIn_0_79, KeyWire_0[79]);
  not KeyNOTGate_0_36(N427, KeyNOTWire_0[36]);
  and AND3_114 (KeyWire_0[80], N393, N17, N287);
  xor KeyGate_0_80(KeyNOTWire_0[37], keyIn_0_80, KeyWire_0[80]);
  not KeyNOTGate_0_37(N432, KeyNOTWire_0[37]);
  nand NAND3_115 (KeyWire_0[81], N393, N287, N55);
  xor KeyGate_0_81(N437, keyIn_0_81, KeyWire_0[81]);
  nand NAND4_116 (KeyWire_0[82], N375, N59, N156, N393);
  xor KeyGate_0_82(N442, keyIn_0_82, KeyWire_0[82]);
  nand NAND3_117 (KeyWire_0[83], N393, N319, N17);
  xor KeyGate_0_83(KeyNOTWire_0[38], keyIn_0_83, KeyWire_0[83]);
  not KeyNOTGate_0_38(N443, KeyNOTWire_0[38]);
  and AND2_118 (KeyWire_0[84], N411, N412);
  xnor KeyGate_0_84(KeyNOTWire_0[39], keyIn_0_84, KeyWire_0[84]);
  not KeyNOTGate_0_39(N444, KeyNOTWire_0[39]);
  and AND2_119 (KeyWire_0[85], N414, N415);
  xnor KeyGate_0_85(KeyNOTWire_0[40], keyIn_0_85, KeyWire_0[85]);
  not KeyNOTGate_0_40(N445, KeyNOTWire_0[40]);
buf BUFF1_120 (N446, N392);
buf BUFF1_121 (N447, N399);
buf BUFF1_122 (N448, N401);
buf BUFF1_123 (N449, N402);
buf BUFF1_124 (N450, N403);
not NOT1_125 (N451, N424);
  nor NOR2_126 (KeyWire_0[86], N406, N425);
  xnor KeyGate_0_86(N460, keyIn_0_86, KeyWire_0[86]);
  nor NOR2_127 (KeyWire_0[87], N409, N426);
  xor KeyGate_0_87(N463, keyIn_0_87, KeyWire_0[87]);
  nand NAND2_128 (KeyWire_0[88], N442, N410);
  xnor KeyGate_0_88(N466, keyIn_0_88, KeyWire_0[88]);
  and AND2_129 (KeyWire_0[89], N143, N427);
  xor KeyGate_0_89(N475, keyIn_0_89, KeyWire_0[89]);
  and AND2_130 (KeyWire_0[90], N310, N432);
  xnor KeyGate_0_90(N476, keyIn_0_90, KeyWire_0[90]);
  and AND2_131 (KeyWire_0[91], N146, N427);
  xor KeyGate_0_91(KeyNOTWire_0[41], keyIn_0_91, KeyWire_0[91]);
  not KeyNOTGate_0_41(N477, KeyNOTWire_0[41]);
  and AND2_132 (KeyWire_0[92], N310, N432);
  xnor KeyGate_0_92(KeyNOTWire_0[42], keyIn_0_92, KeyWire_0[92]);
  not KeyNOTGate_0_42(N478, KeyNOTWire_0[42]);
  and AND2_133 (KeyWire_0[93], N149, N427);
  xor KeyGate_0_93(KeyNOTWire_0[43], keyIn_0_93, KeyWire_0[93]);
  not KeyNOTGate_0_43(N479, KeyNOTWire_0[43]);
  and AND2_134 (KeyWire_0[94], N310, N432);
  xor KeyGate_0_94(N480, keyIn_0_94, KeyWire_0[94]);
  and AND2_135 (KeyWire_0[95], N153, N427);
  xnor KeyGate_0_95(N481, keyIn_0_95, KeyWire_0[95]);
  and AND2_136 (KeyWire_0[96], N310, N432);
  xnor KeyGate_0_96(N482, keyIn_0_96, KeyWire_0[96]);
  nand NAND2_137 (KeyWire_0[97], N443, N1);
  xnor KeyGate_0_97(KeyNOTWire_0[44], keyIn_0_97, KeyWire_0[97]);
  not KeyNOTGate_0_44(N483, KeyNOTWire_0[44]);
  or OR2_138 (KeyWire_0[98], N369, N437);
  xor KeyGate_0_98(N488, keyIn_0_98, KeyWire_0[98]);
  or OR2_139 (KeyWire_0[99], N369, N437);
  xnor KeyGate_0_99(KeyNOTWire_0[45], keyIn_0_99, KeyWire_0[99]);
  not KeyNOTGate_0_45(N489, KeyNOTWire_0[45]);
  or OR2_140 (KeyWire_0[100], N369, N437);
  xor KeyGate_0_100(KeyNOTWire_0[46], keyIn_0_100, KeyWire_0[100]);
  not KeyNOTGate_0_46(N490, KeyNOTWire_0[46]);
or OR2_141 (N491, N369, N437);
  nor NOR2_142 (KeyWire_0[101], N413, N444);
  xnor KeyGate_0_101(KeyNOTWire_0[47], keyIn_0_101, KeyWire_0[101]);
  not KeyNOTGate_0_47(N492, KeyNOTWire_0[47]);
nor NOR2_143 (N495, N416, N445);
  nand NAND2_144 (KeyWire_0[102], N130, N460);
  xor KeyGate_0_102(N498, keyIn_0_102, KeyWire_0[102]);
  or OR2_145 (KeyWire_0[103], N130, N460);
  xnor KeyGate_0_103(N499, keyIn_0_103, KeyWire_0[103]);
  nand NAND2_146 (KeyWire_0[104], N463, N135);
  xor KeyGate_0_104(N500, keyIn_0_104, KeyWire_0[104]);
  or OR2_147 (KeyWire_0[105], N463, N135);
  xnor KeyGate_0_105(N501, keyIn_0_105, KeyWire_0[105]);
and AND2_148 (N502, N91, N466);
nor NOR2_149 (N503, N475, N476);
  and AND2_150 (KeyWire_0[106], N96, N466);
  xor KeyGate_0_106(N504, keyIn_0_106, KeyWire_0[106]);
  nor NOR2_151 (KeyWire_0[107], N477, N478);
  xor KeyGate_0_107(N505, keyIn_0_107, KeyWire_0[107]);
and AND2_152 (N506, N101, N466);
  nor NOR2_153 (KeyWire_0[108], N479, N480);
  xnor KeyGate_0_108(N507, keyIn_0_108, KeyWire_0[108]);
  and AND2_154 (KeyWire_0[109], N106, N466);
  xnor KeyGate_0_109(KeyNOTWire_0[48], keyIn_0_109, KeyWire_0[109]);
  not KeyNOTGate_0_48(N508, KeyNOTWire_0[48]);
  nor NOR2_155 (KeyWire_0[110], N481, N482);
  xor KeyGate_0_110(N509, keyIn_0_110, KeyWire_0[110]);
and AND2_156 (N510, N143, N483);
  and AND2_157 (KeyWire_0[111], N111, N466);
  xnor KeyGate_0_111(N511, keyIn_0_111, KeyWire_0[111]);
and AND2_158 (N512, N146, N483);
and AND2_159 (N513, N116, N466);
  and AND2_160 (KeyWire_0[112], N149, N483);
  xor KeyGate_0_112(KeyNOTWire_0[49], keyIn_0_112, KeyWire_0[112]);
  not KeyNOTGate_0_49(N514, KeyNOTWire_0[49]);
  and AND2_161 (KeyWire_0[113], N121, N466);
  xor KeyGate_0_113(N515, keyIn_0_113, KeyWire_0[113]);
and AND2_162 (N516, N153, N483);
and AND2_163 (N517, N126, N466);
  nand NAND2_164 (KeyWire_0[114], N130, N492);
  xnor KeyGate_0_114(N518, keyIn_0_114, KeyWire_0[114]);
  or OR2_165 (KeyWire_0[115], N130, N492);
  xor KeyGate_0_115(N519, keyIn_0_115, KeyWire_0[115]);
  nand NAND2_166 (KeyWire_0[116], N495, N207);
  xor KeyGate_0_116(N520, keyIn_0_116, KeyWire_0[116]);
or OR2_167 (N521, N495, N207);
  and AND2_168 (KeyWire_0[117], N451, N159);
  xor KeyGate_0_117(KeyNOTWire_0[50], keyIn_0_117, KeyWire_0[117]);
  not KeyNOTGate_0_50(N522, KeyNOTWire_0[50]);
  and AND2_169 (KeyWire_0[118], N451, N165);
  xor KeyGate_0_118(KeyNOTWire_0[51], keyIn_0_118, KeyWire_0[118]);
  not KeyNOTGate_0_51(N523, KeyNOTWire_0[51]);
  and AND2_170 (KeyWire_0[119], N451, N171);
  xor KeyGate_0_119(KeyNOTWire_0[52], keyIn_0_119, KeyWire_0[119]);
  not KeyNOTGate_0_52(N524, KeyNOTWire_0[52]);
  and AND2_171 (KeyWire_0[120], N451, N177);
  xnor KeyGate_0_120(N525, keyIn_0_120, KeyWire_0[120]);
  and AND2_172 (KeyWire_0[121], N451, N183);
  xor KeyGate_0_121(KeyNOTWire_0[53], keyIn_0_121, KeyWire_0[121]);
  not KeyNOTGate_0_53(N526, KeyNOTWire_0[53]);
nand NAND2_173 (N527, N451, N189);
nand NAND2_174 (N528, N451, N195);
nand NAND2_175 (N529, N451, N201);
  nand NAND2_176 (KeyWire_0[122], N498, N499);
  xor KeyGate_0_122(KeyNOTWire_0[54], keyIn_0_122, KeyWire_0[122]);
  not KeyNOTGate_0_54(N530, KeyNOTWire_0[54]);
  nand NAND2_177 (KeyWire_0[123], N500, N501);
  xor KeyGate_0_123(KeyNOTWire_0[55], keyIn_0_123, KeyWire_0[123]);
  not KeyNOTGate_0_55(N533, KeyNOTWire_0[55]);
nor NOR2_178 (N536, N309, N502);
nor NOR2_179 (N537, N316, N504);
  nor NOR2_180 (KeyWire_0[124], N317, N506);
  xor KeyGate_0_124(N538, keyIn_0_124, KeyWire_0[124]);
  nor NOR2_181 (KeyWire_0[125], N318, N508);
  xor KeyGate_0_125(N539, keyIn_0_125, KeyWire_0[125]);
  nor NOR2_182 (KeyWire_0[126], N510, N511);
  xor KeyGate_0_126(N540, keyIn_0_126, KeyWire_0[126]);
nor NOR2_183 (N541, N512, N513);
nor NOR2_184 (N542, N514, N515);
  nor NOR2_185 (KeyWire_0[127], N516, N517);
  xnor KeyGate_0_127(KeyNOTWire_0[56], keyIn_0_127, KeyWire_0[127]);
  not KeyNOTGate_0_56(N543, KeyNOTWire_0[56]);
nand NAND2_186 (N544, N518, N519);
nand NAND2_187 (N547, N520, N521);
  not NOT1_188 (KeyWire_0[128], N530);
  xnor KeyGate_0_128(KeyNOTWire_0[57], keyIn_0_128, KeyWire_0[128]);
  not KeyNOTGate_0_57(N550, KeyNOTWire_0[57]);
  not NOT1_189 (KeyWire_0[129], N533);
  xor KeyGate_0_129(N551, keyIn_0_129, KeyWire_0[129]);
and AND2_190 (N552, N530, N533);
nand NAND2_191 (N553, N536, N503);
  nand NAND2_192 (KeyWire_0[130], N537, N505);
  xor KeyGate_0_130(KeyNOTWire_0[58], keyIn_0_130, KeyWire_0[130]);
  not KeyNOTGate_0_58(N557, KeyNOTWire_0[58]);
  nand NAND2_193 (KeyWire_0[131], N538, N507);
  xnor KeyGate_0_131(KeyNOTWire_0[59], keyIn_0_131, KeyWire_0[131]);
  not KeyNOTGate_0_59(N561, KeyNOTWire_0[59]);
nand NAND2_194 (N565, N539, N509);
  nand NAND2_195 (KeyWire_0[132], N488, N540);
  xor KeyGate_0_132(N569, keyIn_0_132, KeyWire_0[132]);
  nand NAND2_196 (KeyWire_0[133], N489, N541);
  xor KeyGate_0_133(N573, keyIn_0_133, KeyWire_0[133]);
  nand NAND2_197 (KeyWire_0[134], N490, N542);
  xor KeyGate_0_134(KeyNOTWire_0[60], keyIn_0_134, KeyWire_0[134]);
  not KeyNOTGate_0_60(N577, KeyNOTWire_0[60]);
  nand NAND2_198 (KeyWire_0[135], N491, N543);
  xor KeyGate_0_135(N581, keyIn_0_135, KeyWire_0[135]);
  not NOT1_199 (KeyWire_0[136], N544);
  xnor KeyGate_0_136(N585, keyIn_0_136, KeyWire_0[136]);
not NOT1_200 (N586, N547);
  and AND2_201 (KeyWire_0[137], N544, N547);
  xnor KeyGate_0_137(N587, keyIn_0_137, KeyWire_0[137]);
  and AND2_202 (KeyWire_0[138], N550, N551);
  xor KeyGate_0_138(KeyNOTWire_0[61], keyIn_0_138, KeyWire_0[138]);
  not KeyNOTGate_0_61(N588, KeyNOTWire_0[61]);
  and AND2_203 (KeyWire_0[139], N585, N586);
  xnor KeyGate_0_139(KeyNOTWire_0[62], keyIn_0_139, KeyWire_0[139]);
  not KeyNOTGate_0_62(N589, KeyNOTWire_0[62]);
  nand NAND2_204 (KeyWire_0[140], N553, N159);
  xnor KeyGate_0_140(KeyNOTWire_0[63], keyIn_0_140, KeyWire_0[140]);
  not KeyNOTGate_0_63(N590, KeyNOTWire_0[63]);
  or OR2_205 (KeyWire_0[141], N553, N159);
  xnor KeyGate_0_141(KeyNOTWire_0[64], keyIn_0_141, KeyWire_0[141]);
  not KeyNOTGate_0_64(N593, KeyNOTWire_0[64]);
  and AND2_206 (KeyWire_0[142], N246, N553);
  xor KeyGate_0_142(KeyNOTWire_0[65], keyIn_0_142, KeyWire_0[142]);
  not KeyNOTGate_0_65(N596, KeyNOTWire_0[65]);
  nand NAND2_207 (KeyWire_0[143], N557, N165);
  xor KeyGate_0_143(N597, keyIn_0_143, KeyWire_0[143]);
  or OR2_208 (KeyWire_0[144], N557, N165);
  xnor KeyGate_0_144(KeyNOTWire_0[66], keyIn_0_144, KeyWire_0[144]);
  not KeyNOTGate_0_66(N600, KeyNOTWire_0[66]);
and AND2_209 (N605, N246, N557);
nand NAND2_210 (N606, N561, N171);
  or OR2_211 (KeyWire_0[145], N561, N171);
  xnor KeyGate_0_145(N609, keyIn_0_145, KeyWire_0[145]);
and AND2_212 (N615, N246, N561);
  nand NAND2_213 (KeyWire_0[146], N565, N177);
  xor KeyGate_0_146(KeyNOTWire_0[67], keyIn_0_146, KeyWire_0[146]);
  not KeyNOTGate_0_67(N616, KeyNOTWire_0[67]);
  or OR2_214 (KeyWire_0[147], N565, N177);
  xnor KeyGate_0_147(N619, keyIn_0_147, KeyWire_0[147]);
  and AND2_215 (KeyWire_0[148], N246, N565);
  xor KeyGate_0_148(KeyNOTWire_0[68], keyIn_0_148, KeyWire_0[148]);
  not KeyNOTGate_0_68(N624, KeyNOTWire_0[68]);
  nand NAND2_216 (KeyWire_0[149], N569, N183);
  xnor KeyGate_0_149(KeyNOTWire_0[69], keyIn_0_149, KeyWire_0[149]);
  not KeyNOTGate_0_69(N625, KeyNOTWire_0[69]);
  or OR2_217 (KeyWire_0[150], N569, N183);
  xnor KeyGate_0_150(N628, keyIn_0_150, KeyWire_0[150]);
and AND2_218 (N631, N246, N569);
nand NAND2_219 (N632, N573, N189);
or OR2_220 (N635, N573, N189);
  and AND2_221 (KeyWire_0[151], N246, N573);
  xor KeyGate_0_151(KeyNOTWire_0[70], keyIn_0_151, KeyWire_0[151]);
  not KeyNOTGate_0_70(N640, KeyNOTWire_0[70]);
nand NAND2_222 (N641, N577, N195);
  or OR2_223 (KeyWire_0[152], N577, N195);
  xnor KeyGate_0_152(N644, keyIn_0_152, KeyWire_0[152]);
  and AND2_224 (KeyWire_0[153], N246, N577);
  xor KeyGate_0_153(KeyNOTWire_0[71], keyIn_0_153, KeyWire_0[153]);
  not KeyNOTGate_0_71(N650, KeyNOTWire_0[71]);
nand NAND2_225 (N651, N581, N201);
  or OR2_226 (KeyWire_0[154], N581, N201);
  xor KeyGate_0_154(N654, keyIn_0_154, KeyWire_0[154]);
  and AND2_227 (KeyWire_0[155], N246, N581);
  xnor KeyGate_0_155(N659, keyIn_0_155, KeyWire_0[155]);
  nor NOR2_228 (KeyWire_0[156], N552, N588);
  xnor KeyGate_0_156(N660, keyIn_0_156, KeyWire_0[156]);
  nor NOR2_229 (KeyWire_0[157], N587, N589);
  xnor KeyGate_0_157(N661, keyIn_0_157, KeyWire_0[157]);
not NOT1_230 (N662, N590);
  and AND2_231 (KeyWire_0[158], N593, N590);
  xnor KeyGate_0_158(N665, keyIn_0_158, KeyWire_0[158]);
nor NOR2_232 (N669, N596, N522);
not NOT1_233 (N670, N597);
  and AND2_234 (KeyWire_0[159], N600, N597);
  xor KeyGate_0_159(N673, keyIn_0_159, KeyWire_0[159]);
nor NOR2_235 (N677, N605, N523);
not NOT1_236 (N678, N606);
  and AND2_237 (KeyWire_0[160], N609, N606);
  xnor KeyGate_0_160(N682, keyIn_0_160, KeyWire_0[160]);
  nor NOR2_238 (KeyWire_0[161], N615, N524);
  xnor KeyGate_0_161(KeyNOTWire_0[72], keyIn_0_161, KeyWire_0[161]);
  not KeyNOTGate_0_72(N686, KeyNOTWire_0[72]);
  not NOT1_239 (KeyWire_0[162], N616);
  xnor KeyGate_0_162(KeyNOTWire_0[73], keyIn_0_162, KeyWire_0[162]);
  not KeyNOTGate_0_73(N687, KeyNOTWire_0[73]);
  and AND2_240 (KeyWire_0[163], N619, N616);
  xor KeyGate_0_163(KeyNOTWire_0[74], keyIn_0_163, KeyWire_0[163]);
  not KeyNOTGate_0_74(N692, KeyNOTWire_0[74]);
  nor NOR2_241 (KeyWire_0[164], N624, N525);
  xnor KeyGate_0_164(KeyNOTWire_0[75], keyIn_0_164, KeyWire_0[164]);
  not KeyNOTGate_0_75(N696, KeyNOTWire_0[75]);
not NOT1_242 (N697, N625);
  and AND2_243 (KeyWire_0[165], N628, N625);
  xnor KeyGate_0_165(KeyNOTWire_0[76], keyIn_0_165, KeyWire_0[165]);
  not KeyNOTGate_0_76(N700, KeyNOTWire_0[76]);
  nor NOR2_244 (KeyWire_0[166], N631, N526);
  xnor KeyGate_0_166(KeyNOTWire_0[77], keyIn_0_166, KeyWire_0[166]);
  not KeyNOTGate_0_77(N704, KeyNOTWire_0[77]);
not NOT1_245 (N705, N632);
  and AND2_246 (KeyWire_0[167], N635, N632);
  xor KeyGate_0_167(N708, keyIn_0_167, KeyWire_0[167]);
  nor NOR2_247 (KeyWire_0[168], N337, N640);
  xor KeyGate_0_168(N712, keyIn_0_168, KeyWire_0[168]);
  not NOT1_248 (KeyWire_0[169], N641);
  xor KeyGate_0_169(KeyNOTWire_0[78], keyIn_0_169, KeyWire_0[169]);
  not KeyNOTGate_0_78(N713, KeyNOTWire_0[78]);
  and AND2_249 (KeyWire_0[170], N644, N641);
  xor KeyGate_0_170(N717, keyIn_0_170, KeyWire_0[170]);
  nor NOR2_250 (KeyWire_0[171], N339, N650);
  xnor KeyGate_0_171(N721, keyIn_0_171, KeyWire_0[171]);
  not NOT1_251 (KeyWire_0[172], N651);
  xnor KeyGate_0_172(KeyNOTWire_0[79], keyIn_0_172, KeyWire_0[172]);
  not KeyNOTGate_0_79(N722, KeyNOTWire_0[79]);
and AND2_252 (N727, N654, N651);
  nor NOR2_253 (KeyWire_0[173], N341, N659);
  xnor KeyGate_0_173(N731, keyIn_0_173, KeyWire_0[173]);
  nand NAND2_254 (KeyWire_0[174], N654, N261);
  xor KeyGate_0_174(N732, keyIn_0_174, KeyWire_0[174]);
  nand NAND3_255 (KeyWire_0[175], N644, N654, N261);
  xor KeyGate_0_175(KeyNOTWire_0[80], keyIn_0_175, KeyWire_0[175]);
  not KeyNOTGate_0_80(N733, KeyNOTWire_0[80]);
  nand NAND4_256 (KeyWire_0[176], N635, N644, N654, N261);
  xnor KeyGate_0_176(KeyNOTWire_0[81], keyIn_0_176, KeyWire_0[176]);
  not KeyNOTGate_0_81(N734, KeyNOTWire_0[81]);
  not NOT1_257 (KeyWire_0[177], N662);
  xnor KeyGate_0_177(N735, keyIn_0_177, KeyWire_0[177]);
  and AND2_258 (KeyWire_0[178], N228, N665);
  xnor KeyGate_0_178(KeyNOTWire_0[82], keyIn_0_178, KeyWire_0[178]);
  not KeyNOTGate_0_82(N736, KeyNOTWire_0[82]);
and AND2_259 (N737, N237, N662);
  not NOT1_260 (KeyWire_0[179], N670);
  xnor KeyGate_0_179(KeyNOTWire_0[83], keyIn_0_179, KeyWire_0[179]);
  not KeyNOTGate_0_83(N738, KeyNOTWire_0[83]);
  and AND2_261 (KeyWire_0[180], N228, N673);
  xnor KeyGate_0_180(N739, keyIn_0_180, KeyWire_0[180]);
and AND2_262 (N740, N237, N670);
  not NOT1_263 (KeyWire_0[181], N678);
  xnor KeyGate_0_181(N741, keyIn_0_181, KeyWire_0[181]);
and AND2_264 (N742, N228, N682);
  and AND2_265 (KeyWire_0[182], N237, N678);
  xnor KeyGate_0_182(N743, keyIn_0_182, KeyWire_0[182]);
  not NOT1_266 (KeyWire_0[183], N687);
  xnor KeyGate_0_183(KeyNOTWire_0[84], keyIn_0_183, KeyWire_0[183]);
  not KeyNOTGate_0_84(N744, KeyNOTWire_0[84]);
  and AND2_267 (KeyWire_0[184], N228, N692);
  xor KeyGate_0_184(KeyNOTWire_0[85], keyIn_0_184, KeyWire_0[184]);
  not KeyNOTGate_0_85(N745, KeyNOTWire_0[85]);
and AND2_268 (N746, N237, N687);
  not NOT1_269 (KeyWire_0[185], N697);
  xor KeyGate_0_185(N747, keyIn_0_185, KeyWire_0[185]);
and AND2_270 (N748, N228, N700);
  and AND2_271 (KeyWire_0[186], N237, N697);
  xor KeyGate_0_186(KeyNOTWire_0[86], keyIn_0_186, KeyWire_0[186]);
  not KeyNOTGate_0_86(N749, KeyNOTWire_0[86]);
not NOT1_272 (N750, N705);
  and AND2_273 (KeyWire_0[187], N228, N708);
  xor KeyGate_0_187(KeyNOTWire_0[87], keyIn_0_187, KeyWire_0[187]);
  not KeyNOTGate_0_87(N751, KeyNOTWire_0[87]);
  and AND2_274 (KeyWire_0[188], N237, N705);
  xnor KeyGate_0_188(N752, keyIn_0_188, KeyWire_0[188]);
  not NOT1_275 (KeyWire_0[189], N713);
  xor KeyGate_0_189(KeyNOTWire_0[88], keyIn_0_189, KeyWire_0[189]);
  not KeyNOTGate_0_88(N753, KeyNOTWire_0[88]);
  and AND2_276 (KeyWire_0[190], N228, N717);
  xor KeyGate_0_190(N754, keyIn_0_190, KeyWire_0[190]);
  and AND2_277 (KeyWire_0[191], N237, N713);
  xor KeyGate_0_191(KeyNOTWire_0[89], keyIn_0_191, KeyWire_0[191]);
  not KeyNOTGate_0_89(N755, KeyNOTWire_0[89]);
not NOT1_278 (N756, N722);
nor NOR2_279 (N757, N727, N261);
  and AND2_280 (KeyWire_0[192], N727, N261);
  xnor KeyGate_0_192(KeyNOTWire_0[90], keyIn_0_192, KeyWire_0[192]);
  not KeyNOTGate_0_90(N758, KeyNOTWire_0[90]);
  and AND2_281 (KeyWire_0[193], N228, N727);
  xnor KeyGate_0_193(KeyNOTWire_0[91], keyIn_0_193, KeyWire_0[193]);
  not KeyNOTGate_0_91(N759, KeyNOTWire_0[91]);
  and AND2_282 (KeyWire_0[194], N237, N722);
  xnor KeyGate_0_194(N760, keyIn_0_194, KeyWire_0[194]);
  nand NAND2_283 (KeyWire_0[195], N644, N722);
  xnor KeyGate_0_195(N761, keyIn_0_195, KeyWire_0[195]);
  nand NAND2_284 (KeyWire_0[196], N635, N713);
  xnor KeyGate_0_196(N762, keyIn_0_196, KeyWire_0[196]);
  nand NAND3_285 (KeyWire_0[197], N635, N644, N722);
  xnor KeyGate_0_197(KeyNOTWire_0[92], keyIn_0_197, KeyWire_0[197]);
  not KeyNOTGate_0_92(N763, KeyNOTWire_0[92]);
  nand NAND2_286 (KeyWire_0[198], N609, N687);
  xor KeyGate_0_198(N764, keyIn_0_198, KeyWire_0[198]);
  nand NAND2_287 (KeyWire_0[199], N600, N678);
  xnor KeyGate_0_199(KeyNOTWire_0[93], keyIn_0_199, KeyWire_0[199]);
  not KeyNOTGate_0_93(N765, KeyNOTWire_0[93]);
  nand NAND3_288 (KeyWire_0[200], N600, N609, N687);
  xnor KeyGate_0_200(KeyNOTWire_0[94], keyIn_0_200, KeyWire_0[200]);
  not KeyNOTGate_0_94(N766, KeyNOTWire_0[94]);
buf BUFF1_289 (N767, N660);
buf BUFF1_290 (N768, N661);
  nor NOR2_291 (KeyWire_0[201], N736, N737);
  xor KeyGate_0_201(N769, keyIn_0_201, KeyWire_0[201]);
  nor NOR2_292 (KeyWire_0[202], N739, N740);
  xor KeyGate_0_202(N770, keyIn_0_202, KeyWire_0[202]);
  nor NOR2_293 (KeyWire_0[203], N742, N743);
  xnor KeyGate_0_203(KeyNOTWire_0[95], keyIn_0_203, KeyWire_0[203]);
  not KeyNOTGate_0_95(N771, KeyNOTWire_0[95]);
nor NOR2_294 (N772, N745, N746);
  nand NAND4_295 (KeyWire_0[204], N750, N762, N763, N734);
  xor KeyGate_0_204(N773, keyIn_0_204, KeyWire_0[204]);
  nor NOR2_296 (KeyWire_0[205], N748, N749);
  xnor KeyGate_0_205(N777, keyIn_0_205, KeyWire_0[205]);
  nand NAND3_297 (KeyWire_0[206], N753, N761, N733);
  xor KeyGate_0_206(KeyNOTWire_0[96], keyIn_0_206, KeyWire_0[206]);
  not KeyNOTGate_0_96(N778, KeyNOTWire_0[96]);
nor NOR2_298 (N781, N751, N752);
  nand NAND2_299 (KeyWire_0[207], N756, N732);
  xor KeyGate_0_207(N782, keyIn_0_207, KeyWire_0[207]);
  nor NOR2_300 (KeyWire_0[208], N754, N755);
  xor KeyGate_0_208(N785, keyIn_0_208, KeyWire_0[208]);
  nor NOR2_301 (KeyWire_0[209], N757, N758);
  xor KeyGate_0_209(KeyNOTWire_0[97], keyIn_0_209, KeyWire_0[209]);
  not KeyNOTGate_0_97(N786, KeyNOTWire_0[97]);
  nor NOR2_302 (KeyWire_0[210], N759, N760);
  xor KeyGate_0_210(N787, keyIn_0_210, KeyWire_0[210]);
  nor NOR2_303 (KeyWire_0[211], N700, N773);
  xnor KeyGate_0_211(N788, keyIn_0_211, KeyWire_0[211]);
and AND2_304 (N789, N700, N773);
nor NOR2_305 (N790, N708, N778);
  and AND2_306 (KeyWire_0[212], N708, N778);
  xor KeyGate_0_212(KeyNOTWire_0[98], keyIn_0_212, KeyWire_0[212]);
  not KeyNOTGate_0_98(N791, KeyNOTWire_0[98]);
  nor NOR2_307 (KeyWire_0[213], N717, N782);
  xnor KeyGate_0_213(KeyNOTWire_0[99], keyIn_0_213, KeyWire_0[213]);
  not KeyNOTGate_0_99(N792, KeyNOTWire_0[99]);
  and AND2_308 (KeyWire_0[214], N717, N782);
  xnor KeyGate_0_214(KeyNOTWire_0[100], keyIn_0_214, KeyWire_0[214]);
  not KeyNOTGate_0_100(N793, KeyNOTWire_0[100]);
  and AND2_309 (KeyWire_0[215], N219, N786);
  xor KeyGate_0_215(N794, keyIn_0_215, KeyWire_0[215]);
nand NAND2_310 (N795, N628, N773);
nand NAND2_311 (N796, N795, N747);
  nor NOR2_312 (KeyWire_0[216], N788, N789);
  xor KeyGate_0_216(KeyNOTWire_0[101], keyIn_0_216, KeyWire_0[216]);
  not KeyNOTGate_0_101(N802, KeyNOTWire_0[101]);
nor NOR2_313 (N803, N790, N791);
  nor NOR2_314 (KeyWire_0[217], N792, N793);
  xnor KeyGate_0_217(KeyNOTWire_0[102], keyIn_0_217, KeyWire_0[217]);
  not KeyNOTGate_0_102(N804, KeyNOTWire_0[102]);
nor NOR2_315 (N805, N340, N794);
  nor NOR2_316 (KeyWire_0[218], N692, N796);
  xnor KeyGate_0_218(N806, keyIn_0_218, KeyWire_0[218]);
  and AND2_317 (KeyWire_0[219], N692, N796);
  xnor KeyGate_0_219(KeyNOTWire_0[103], keyIn_0_219, KeyWire_0[219]);
  not KeyNOTGate_0_103(N807, KeyNOTWire_0[103]);
  and AND2_318 (KeyWire_0[220], N219, N802);
  xnor KeyGate_0_220(KeyNOTWire_0[104], keyIn_0_220, KeyWire_0[220]);
  not KeyNOTGate_0_104(N808, KeyNOTWire_0[104]);
  and AND2_319 (KeyWire_0[221], N219, N803);
  xnor KeyGate_0_221(N809, keyIn_0_221, KeyWire_0[221]);
  and AND2_320 (KeyWire_0[222], N219, N804);
  xor KeyGate_0_222(KeyNOTWire_0[105], keyIn_0_222, KeyWire_0[222]);
  not KeyNOTGate_0_105(N810, KeyNOTWire_0[105]);
  nand NAND4_321 (KeyWire_0[223], N805, N787, N731, N529);
  xnor KeyGate_0_223(KeyNOTWire_0[106], keyIn_0_223, KeyWire_0[223]);
  not KeyNOTGate_0_106(N811, KeyNOTWire_0[106]);
nand NAND2_322 (N812, N619, N796);
  nand NAND3_323 (KeyWire_0[224], N609, N619, N796);
  xor KeyGate_0_224(KeyNOTWire_0[107], keyIn_0_224, KeyWire_0[224]);
  not KeyNOTGate_0_107(N813, KeyNOTWire_0[107]);
  nand NAND4_324 (KeyWire_0[225], N600, N609, N619, N796);
  xor KeyGate_0_225(N814, keyIn_0_225, KeyWire_0[225]);
nand NAND4_325 (N815, N738, N765, N766, N814);
nand NAND3_326 (N819, N741, N764, N813);
nand NAND2_327 (N822, N744, N812);
nor NOR2_328 (N825, N806, N807);
  nor NOR2_329 (KeyWire_0[226], N335, N808);
  xor KeyGate_0_226(KeyNOTWire_0[108], keyIn_0_226, KeyWire_0[226]);
  not KeyNOTGate_0_108(N826, KeyNOTWire_0[108]);
  nor NOR2_330 (KeyWire_0[227], N336, N809);
  xor KeyGate_0_227(N827, keyIn_0_227, KeyWire_0[227]);
  nor NOR2_331 (KeyWire_0[228], N338, N810);
  xnor KeyGate_0_228(KeyNOTWire_0[109], keyIn_0_228, KeyWire_0[228]);
  not KeyNOTGate_0_109(N828, KeyNOTWire_0[109]);
  not NOT1_332 (KeyWire_0[229], N811);
  xor KeyGate_0_229(N829, keyIn_0_229, KeyWire_0[229]);
nor NOR2_333 (N830, N665, N815);
  and AND2_334 (KeyWire_0[230], N665, N815);
  xor KeyGate_0_230(KeyNOTWire_0[110], keyIn_0_230, KeyWire_0[230]);
  not KeyNOTGate_0_110(N831, KeyNOTWire_0[110]);
nor NOR2_335 (N832, N673, N819);
and AND2_336 (N833, N673, N819);
  nor NOR2_337 (KeyWire_0[231], N682, N822);
  xor KeyGate_0_231(KeyNOTWire_0[111], keyIn_0_231, KeyWire_0[231]);
  not KeyNOTGate_0_111(N834, KeyNOTWire_0[111]);
  and AND2_338 (KeyWire_0[232], N682, N822);
  xnor KeyGate_0_232(KeyNOTWire_0[112], keyIn_0_232, KeyWire_0[232]);
  not KeyNOTGate_0_112(N835, KeyNOTWire_0[112]);
and AND2_339 (N836, N219, N825);
  nand NAND3_340 (KeyWire_0[233], N826, N777, N704);
  xnor KeyGate_0_233(N837, keyIn_0_233, KeyWire_0[233]);
nand NAND4_341 (N838, N827, N781, N712, N527);
nand NAND4_342 (N839, N828, N785, N721, N528);
  not NOT1_343 (KeyWire_0[234], N829);
  xnor KeyGate_0_234(N840, keyIn_0_234, KeyWire_0[234]);
  nand NAND2_344 (KeyWire_0[235], N815, N593);
  xor KeyGate_0_235(KeyNOTWire_0[113], keyIn_0_235, KeyWire_0[235]);
  not KeyNOTGate_0_113(N841, KeyNOTWire_0[113]);
  nor NOR2_345 (KeyWire_0[236], N830, N831);
  xor KeyGate_0_236(KeyNOTWire_0[114], keyIn_0_236, KeyWire_0[236]);
  not KeyNOTGate_0_114(N842, KeyNOTWire_0[114]);
nor NOR2_346 (N843, N832, N833);
  nor NOR2_347 (KeyWire_0[237], N834, N835);
  xnor KeyGate_0_237(KeyNOTWire_0[115], keyIn_0_237, KeyWire_0[237]);
  not KeyNOTGate_0_115(N844, KeyNOTWire_0[115]);
nor NOR2_348 (N845, N334, N836);
  not NOT1_349 (KeyWire_0[238], N837);
  xnor KeyGate_0_238(KeyNOTWire_0[116], keyIn_0_238, KeyWire_0[238]);
  not KeyNOTGate_0_116(N846, KeyNOTWire_0[116]);
  not NOT1_350 (KeyWire_0[239], N838);
  xor KeyGate_0_239(KeyNOTWire_0[117], keyIn_0_239, KeyWire_0[239]);
  not KeyNOTGate_0_117(N847, KeyNOTWire_0[117]);
  not NOT1_351 (KeyWire_0[240], N839);
  xnor KeyGate_0_240(N848, keyIn_0_240, KeyWire_0[240]);
  and AND2_352 (KeyWire_0[241], N735, N841);
  xor KeyGate_0_241(N849, keyIn_0_241, KeyWire_0[241]);
buf BUFF1_353 (N850, N840);
and AND2_354 (N851, N219, N842);
  and AND2_355 (KeyWire_0[242], N219, N843);
  xor KeyGate_0_242(KeyNOTWire_0[118], keyIn_0_242, KeyWire_0[242]);
  not KeyNOTGate_0_118(N852, KeyNOTWire_0[118]);
  and AND2_356 (KeyWire_0[243], N219, N844);
  xor KeyGate_0_243(N853, keyIn_0_243, KeyWire_0[243]);
  nand NAND3_357 (KeyWire_0[244], N845, N772, N696);
  xor KeyGate_0_244(N854, keyIn_0_244, KeyWire_0[244]);
  not NOT1_358 (KeyWire_0[245], N846);
  xnor KeyGate_0_245(KeyNOTWire_0[119], keyIn_0_245, KeyWire_0[245]);
  not KeyNOTGate_0_119(N855, KeyNOTWire_0[119]);
  not NOT1_359 (KeyWire_0[246], N847);
  xor KeyGate_0_246(N856, keyIn_0_246, KeyWire_0[246]);
  not NOT1_360 (KeyWire_0[247], N848);
  xnor KeyGate_0_247(KeyNOTWire_0[120], keyIn_0_247, KeyWire_0[247]);
  not KeyNOTGate_0_120(N857, KeyNOTWire_0[120]);
  not NOT1_361 (KeyWire_0[248], N849);
  xor KeyGate_0_248(KeyNOTWire_0[121], keyIn_0_248, KeyWire_0[248]);
  not KeyNOTGate_0_121(N858, KeyNOTWire_0[121]);
  nor NOR2_362 (KeyWire_0[249], N417, N851);
  xnor KeyGate_0_249(N859, keyIn_0_249, KeyWire_0[249]);
  nor NOR2_363 (KeyWire_0[250], N332, N852);
  xnor KeyGate_0_250(N860, keyIn_0_250, KeyWire_0[250]);
nor NOR2_364 (N861, N333, N853);
not NOT1_365 (N862, N854);
buf BUFF1_366 (N863, N855);
buf BUFF1_367 (N864, N856);
buf BUFF1_368 (N865, N857);
buf BUFF1_369 (N866, N858);
  nand NAND3_370 (KeyWire_0[251], N859, N769, N669);
  xor KeyGate_0_251(KeyNOTWire_0[122], keyIn_0_251, KeyWire_0[251]);
  not KeyNOTGate_0_122(N867, KeyNOTWire_0[122]);
nand NAND3_371 (N868, N860, N770, N677);
  nand NAND3_372 (KeyWire_0[252], N861, N771, N686);
  xor KeyGate_0_252(KeyNOTWire_0[123], keyIn_0_252, KeyWire_0[252]);
  not KeyNOTGate_0_123(N869, KeyNOTWire_0[123]);
  not NOT1_373 (KeyWire_0[253], N862);
  xnor KeyGate_0_253(KeyNOTWire_0[124], keyIn_0_253, KeyWire_0[253]);
  not KeyNOTGate_0_124(N870, KeyNOTWire_0[124]);
  not NOT1_374 (KeyWire_0[254], N867);
  xnor KeyGate_0_254(KeyNOTWire_0[125], keyIn_0_254, KeyWire_0[254]);
  not KeyNOTGate_0_125(N871, KeyNOTWire_0[125]);
  not NOT1_375 (KeyWire_0[255], N868);
  xor KeyGate_0_255(N872, keyIn_0_255, KeyWire_0[255]);
not NOT1_376 (N873, N869);
buf BUFF1_377 (N874, N870);
not NOT1_378 (N875, N871);
not NOT1_379 (N876, N872);
not NOT1_380 (N877, N873);
buf BUFF1_381 (N878, N875);
buf BUFF1_382 (N879, N876);
buf BUFF1_383 (N880, N877);

endmodule
