`timescale 1ns / 1ps
// Verilog
// c880
// Ninputs 60
// Noutputs 26
// NtotalGates 383
// NAND4 13
// AND3 12
// NAND2 60
// NAND3 14
// AND2 105
// OR2 29
// NOT1 63
// NOR2 61
// BUFF1 26

module top (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
                  N865,N866,N874,N878,N879,N880,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
        keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
                  keyinput125, keyinput126, keyinput127,
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202,
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207,
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212,
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217,
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222,
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227,
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232,
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237,
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242,
                  keyinput243, keyinput244, keyinput245, keyinput246, keyinput247,
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
        keyinput253, keyinput254, keyinput255, keyinput256, keyinput257,
        keyinput258, keyinput259, keyinput260, keyinput261, keyinput262,
        keyinput263, keyinput264, keyinput265, keyinput266, keyinput267,
        keyinput268, keyinput269, keyinput270, keyinput271, keyinput272,
        keyinput273, keyinput274, keyinput275, keyinput276, keyinput277,
        keyinput278, keyinput279, keyinput280, keyinput281, keyinput282,
        keyinput283, keyinput284, keyinput285, keyinput286, keyinput287,
        keyinput288, keyinput289, keyinput290, keyinput291, keyinput292,
        keyinput293, keyinput294, keyinput295, keyinput296, keyinput297,
        keyinput298, keyinput299, keyinput300, keyinput301, keyinput302,
        keyinput303, keyinput304, keyinput305, keyinput306, keyinput307);

  input keyinput248, keyinput249, keyinput250, keyinput251, keyinput252;
  input keyinput253, keyinput254, keyinput255, keyinput256, keyinput257;
  input keyinput258, keyinput259, keyinput260, keyinput261, keyinput262;
  input keyinput263, keyinput264, keyinput265, keyinput266, keyinput267;
  input keyinput268, keyinput269, keyinput270, keyinput271, keyinput272;
  input keyinput273, keyinput274, keyinput275, keyinput276, keyinput277;
  input keyinput278, keyinput279, keyinput280, keyinput281, keyinput282;
  input keyinput283, keyinput284, keyinput285, keyinput286, keyinput287;
  input keyinput288, keyinput289, keyinput290, keyinput291, keyinput292;
  input keyinput293, keyinput294, keyinput295, keyinput296, keyinput297;
  input keyinput298, keyinput299, keyinput300, keyinput301, keyinput302;
  input keyinput303, keyinput304, keyinput305, keyinput306, keyinput307;


  input keyinput128, keyinput129, keyinput130, keyinput131, keyinput132;
  input keyinput133, keyinput134, keyinput135, keyinput136, keyinput137;
  input keyinput138, keyinput139, keyinput140, keyinput141, keyinput142;
  input keyinput143, keyinput144, keyinput145, keyinput146, keyinput147;
  input keyinput148, keyinput149, keyinput150, keyinput151, keyinput152;
  input keyinput153, keyinput154, keyinput155, keyinput156, keyinput157;
  input keyinput158, keyinput159, keyinput160, keyinput161, keyinput162;
  input keyinput163, keyinput164, keyinput165, keyinput166, keyinput167;
  input keyinput168, keyinput169, keyinput170, keyinput171, keyinput172;
  input keyinput173, keyinput174, keyinput175, keyinput176, keyinput177;
  input keyinput178, keyinput179, keyinput180, keyinput181, keyinput182;
  input keyinput183, keyinput184, keyinput185, keyinput186, keyinput187;
  input keyinput188, keyinput189, keyinput190, keyinput191, keyinput192;
  input keyinput193, keyinput194, keyinput195, keyinput196, keyinput197;
  input keyinput198, keyinput199, keyinput200, keyinput201, keyinput202;
  input keyinput203, keyinput204, keyinput205, keyinput206, keyinput207;
  input keyinput208, keyinput209, keyinput210, keyinput211, keyinput212;
  input keyinput213, keyinput214, keyinput215, keyinput216, keyinput217;
  input keyinput218, keyinput219, keyinput220, keyinput221, keyinput222;
  input keyinput223, keyinput224, keyinput225, keyinput226, keyinput227;
  input keyinput228, keyinput229, keyinput230, keyinput231, keyinput232;
  input keyinput233, keyinput234, keyinput235, keyinput236, keyinput237;
  input keyinput238, keyinput239, keyinput240, keyinput241, keyinput242;
  input keyinput243, keyinput244, keyinput245, keyinput246, keyinput247;

  wire KeyWire_0_1 , KeyWire_0_2, keyinput_Wire_1;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31, keyinput32, keyinput33, keyinput34;
  input keyinput35, keyinput36, keyinput37, keyinput38, keyinput39;
  input keyinput40, keyinput41, keyinput42, keyinput43, keyinput44;
  input keyinput45, keyinput46, keyinput47, keyinput48, keyinput49;
  input keyinput50, keyinput51, keyinput52, keyinput53, keyinput54;
  input keyinput55, keyinput56, keyinput57, keyinput58, keyinput59;
  input keyinput60, keyinput61, keyinput62, keyinput63, keyinput64;
  input keyinput65, keyinput66, keyinput67, keyinput68, keyinput69;
  input keyinput70, keyinput71, keyinput72, keyinput73, keyinput74;
  input keyinput75, keyinput76, keyinput77, keyinput78, keyinput79;
  input keyinput80, keyinput81, keyinput82, keyinput83, keyinput84;
  input keyinput85, keyinput86, keyinput87, keyinput88, keyinput89;
  input keyinput90, keyinput91, keyinput92, keyinput93, keyinput94;
  input keyinput95, keyinput96, keyinput97, keyinput98, keyinput99;
  input keyinput100, keyinput101, keyinput102, keyinput103, keyinput104;
  input keyinput105, keyinput106, keyinput107, keyinput108, keyinput109;
  input keyinput110, keyinput111, keyinput112, keyinput113, keyinput114;
  input keyinput115, keyinput116, keyinput117, keyinput118, keyinput119;
  input keyinput120, keyinput121, keyinput122, keyinput123, keyinput124;
  input keyinput125, keyinput126, keyinput127;

  wire [0:127] keyinput_Wire_0;
  wire [0:66] KeyNOTWire_0;

input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;

output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;

wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877;

nand NAND4_1 (N269, N1, N8, N13, N17);
nand NAND4_2 (N270, N1, N26, N13, N17);
and AND3_3 (N273, N29, N36, N42);
  and AND3_4 (keyinput_Wire_0[0], N1, N26, N51);
  xor keyGate_0_0(N276, keyinput0, keyinput_Wire_0[0]);
  nand NAND4_5 (keyinput_Wire_0[1], N1, N8, N51, N17);
  xor keyGate_0_1(N279, keyinput1, keyinput_Wire_0[1]);
nand NAND4_6 (N280, N1, N8, N13, N55);
nand NAND4_7 (N284, N59, N42, N68, N72);
nand NAND2_8 (N285, N29, N68);
nand NAND3_9 (N286, N59, N68, N74);
  and AND3_10 (keyinput_Wire_0[2], N29, N75, N80);
  xnor keyGate_0_2(KeyNOTWire_0[0], keyinput2, keyinput_Wire_0[2]);
  not KeyNOTGate_0_0(N287, KeyNOTWire_0[0]);
and AND3_11 (N290, N29, N75, N42);
and AND3_12 (N291, N29, N36, N80);
and AND3_13 (N292, N29, N36, N42);
and AND3_14 (N293, N59, N75, N80);
  and AND3_15 (keyinput_Wire_0[3], N59, N75, N42);
  xor keyGate_0_3(N294, keyinput3, keyinput_Wire_0[3]);
and AND3_16 (N295, N59, N36, N80);
and AND3_17 (N296, N59, N36, N42);
and AND2_18 (N297, N85, N86);
or OR2_19 (N298, N87, N88);
nand NAND2_20 (N301, N91, N96);
or OR2_21 (N302, N91, N96);
nand NAND2_22 (N303, N101, N106);
or OR2_23 (N304, N101, N106);
nand NAND2_24 (N305, N111, N116);
or OR2_25 (N306, N111, N116);
nand NAND2_26 (N307, N121, N126);
or OR2_27 (N308, N121, N126);
and AND2_28 (N309, N8, N138);
  not NOT1_29 (keyinput_Wire_0[4], N268);
  xnor keyGate_0_4(KeyNOTWire_0[1], keyinput4, keyinput_Wire_0[4]);
  not KeyNOTGate_0_1(N310, KeyNOTWire_0[1]);
and AND2_30 (N316, N51, N138);
and AND2_31 (N317, N17, N138);
and AND2_32 (N318, N152, N138);
  nand NAND2_33 (keyinput_Wire_0[5], N59, N156);
  xor keyGate_0_5(N319, keyinput5, keyinput_Wire_0[5]);
  nor NOR2_34 (keyinput_Wire_0[6], N17, N42);
  xor keyGate_0_6(KeyNOTWire_0[2], keyinput6, keyinput_Wire_0[6]);
  not KeyNOTGate_0_2(N322, KeyNOTWire_0[2]);
  and AND2_35 (keyinput_Wire_0[7], N17, N42);
  xnor keyGate_0_7(KeyNOTWire_0[3], keyinput7, keyinput_Wire_0[7]);
  not KeyNOTGate_0_3(N323, KeyNOTWire_0[3]);
nand NAND2_36 (N324, N159, N165);
or OR2_37 (N325, N159, N165);
nand NAND2_38 (N326, N171, N177);
or OR2_39 (N327, N171, N177);
nand NAND2_40 (N328, N183, N189);
or OR2_41 (N329, N183, N189);
nand NAND2_42 (N330, N195, N201);
or OR2_43 (N331, N195, N201);
and AND2_44 (N332, N210, N91);
and AND2_45 (N333, N210, N96);
and AND2_46 (N334, N210, N101);
and AND2_47 (N335, N210, N106);
and AND2_48 (N336, N210, N111);
and AND2_49 (N337, N255, N259);
and AND2_50 (N338, N210, N116);
and AND2_51 (N339, N255, N260);
and AND2_52 (N340, N210, N121);
and AND2_53 (N341, N255, N267);
not NOT1_54 (N342, N269);
not NOT1_55 (N343, N273);
or OR2_56 (N344, N270, N273);
  not NOT1_57 (keyinput_Wire_0[8], N276);
  xnor keyGate_0_8(N345, keyinput8, keyinput_Wire_0[8]);
not NOT1_58 (N346, N276);
  not NOT1_59 (keyinput_Wire_0[9], N279);
  xor keyGate_0_9(KeyNOTWire_0[4], keyinput9, keyinput_Wire_0[9]);
  not KeyNOTGate_0_4(N347, KeyNOTWire_0[4]);
nor NOR2_60 (N348, N280, N284);
or OR2_61 (N349, N280, N285);
or OR2_62 (N350, N280, N286);
not NOT1_63 (N351, N293);
  not NOT1_64 (keyinput_Wire_0[10], N294);
  xor keyGate_0_10(KeyNOTWire_0[5], keyinput10, keyinput_Wire_0[10]);
  not KeyNOTGate_0_5(N352, KeyNOTWire_0[5]);
not NOT1_65 (N353, N295);
not NOT1_66 (N354, N296);
nand NAND2_67 (N355, N89, N298);
and AND2_68 (N356, N90, N298);
nand NAND2_69 (N357, N301, N302);
nand NAND2_70 (N360, N303, N304);
nand NAND2_71 (N363, N305, N306);
nand NAND2_72 (N366, N307, N308);
  not NOT1_73 (keyinput_Wire_0[11], N310);
  xnor keyGate_0_11(KeyNOTWire_0[6], keyinput11, keyinput_Wire_0[11]);
  not KeyNOTGate_0_6(N369, KeyNOTWire_0[6]);
  nor NOR2_74 (keyinput_Wire_0[12], N322, N323);
  xnor keyGate_0_12(N375, keyinput12, keyinput_Wire_0[12]);
nand NAND2_75 (N376, N324, N325);
nand NAND2_76 (N379, N326, N327);
nand NAND2_77 (N382, N328, N329);
nand NAND2_78 (N385, N330, N331);
buf BUFF1_79 (N388, N290);
buf BUFF1_80 (N389, N291);
buf BUFF1_81 (N390, N292);
buf BUFF1_82 (N391, N297);
or OR2_83 (N392, N270, N343);
  not NOT1_84 (keyinput_Wire_0[13], N345);
  xnor keyGate_0_13(KeyNOTWire_0[7], keyinput13, keyinput_Wire_0[13]);
  not KeyNOTGate_0_7(N393, KeyNOTWire_0[7]);
not NOT1_85 (N399, N346);
and AND2_86 (N400, N348, N73);
not NOT1_87 (N401, N349);
not NOT1_88 (N402, N350);
not NOT1_89 (N403, N355);
not NOT1_90 (N404, N357);
not NOT1_91 (N405, N360);
and AND2_92 (N406, N357, N360);
not NOT1_93 (N407, N363);
not NOT1_94 (N408, N366);
and AND2_95 (N409, N363, N366);
  nand NAND2_96 (keyinput_Wire_0[14], N347, N352);
  xor keyGate_0_14(N410, keyinput14, keyinput_Wire_0[14]);
not NOT1_97 (N411, N376);
not NOT1_98 (N412, N379);
and AND2_99 (N413, N376, N379);
not NOT1_100 (N414, N382);
not NOT1_101 (N415, N385);
and AND2_102 (N416, N382, N385);
and AND2_103 (N417, N210, N369);
buf BUFF1_104 (N418, N342);
buf BUFF1_105 (N419, N344);
buf BUFF1_106 (N420, N351);
buf BUFF1_107 (N421, N353);
buf BUFF1_108 (N422, N354);
buf BUFF1_109 (N423, N356);
not NOT1_110 (N424, N400);
and AND2_111 (N425, N404, N405);
and AND2_112 (N426, N407, N408);
  and AND3_113 (keyinput_Wire_0[15], N319, N393, N55);
  xnor keyGate_0_15(KeyNOTWire_0[8], keyinput15, keyinput_Wire_0[15]);
  not KeyNOTGate_0_8(N427, KeyNOTWire_0[8]);
  and AND3_114 (keyinput_Wire_0[16], N393, N17, N287);
  xor keyGate_0_16(N432, keyinput16, keyinput_Wire_0[16]);
  nand NAND3_115 (keyinput_Wire_0[17], N393, N287, N55);
  xnor keyGate_0_17(N437, keyinput17, keyinput_Wire_0[17]);
  nand NAND4_116 (keyinput_Wire_0[18], N375, N59, N156, N393);
  xnor keyGate_0_18(N442, keyinput18, keyinput_Wire_0[18]);
  nand NAND3_117 (keyinput_Wire_0[19], N393, N319, N17);
  xor keyGate_0_19(KeyNOTWire_0[9], keyinput19, keyinput_Wire_0[19]);
  not KeyNOTGate_0_9(N443, KeyNOTWire_0[9]);
and AND2_118 (N444, N411, N412);
and AND2_119 (N445, N414, N415);
buf BUFF1_120 (N446, N392);
buf BUFF1_121 (N447, N399);
buf BUFF1_122 (N448, N401);
buf BUFF1_123 (N449, N402);
buf BUFF1_124 (N450, N403);
not NOT1_125 (N451, N424);
nor NOR2_126 (N460, N406, N425);
nor NOR2_127 (N463, N409, N426);
  nand NAND2_128 (keyinput_Wire_0[20], N442, N410);
  xor keyGate_0_20(N466, keyinput20, keyinput_Wire_0[20]);
and AND2_129 (N475, N143, N427);
and AND2_130 (N476, N310, N432);
and AND2_131 (N477, N146, N427);
and AND2_132 (N478, N310, N432);
and AND2_133 (N479, N149, N427);
and AND2_134 (N480, N310, N432);
and AND2_135 (N481, N153, N427);
and AND2_136 (N482, N310, N432);
  nand NAND2_137 (keyinput_Wire_0[21], N443, N1);
  xnor keyGate_0_21(N483, keyinput21, keyinput_Wire_0[21]);
or OR2_138 (N488, N369, N437);
  or OR2_139 (keyinput_Wire_0[22], N369, N437);
  xnor keyGate_0_22(N489, keyinput22, keyinput_Wire_0[22]);
  or OR2_140 (keyinput_Wire_0[23], N369, N437);
  xor keyGate_0_23(N490, keyinput23, keyinput_Wire_0[23]);
  or OR2_141 (keyinput_Wire_0[24], N369, N437);
  xor keyGate_0_24(KeyNOTWire_0[10], keyinput24, keyinput_Wire_0[24]);
  not KeyNOTGate_0_10(N491, KeyNOTWire_0[10]);
nor NOR2_142 (N492, N413, N444);
nor NOR2_143 (N495, N416, N445);
nand NAND2_144 (N498, N130, N460);
or OR2_145 (N499, N130, N460);
nand NAND2_146 (N500, N463, N135);
or OR2_147 (N501, N463, N135);
and AND2_148 (N502, N91, N466);
nor NOR2_149 (N503, N475, N476);
and AND2_150 (N504, N96, N466);
nor NOR2_151 (N505, N477, N478);
and AND2_152 (N506, N101, N466);
nor NOR2_153 (N507, N479, N480);
and AND2_154 (N508, N106, N466);
nor NOR2_155 (N509, N481, N482);
and AND2_156 (N510, N143, N483);
  and AND2_157 (keyinput_Wire_0[25], N111, N466);
  xnor keyGate_0_25(N511, keyinput25, keyinput_Wire_0[25]);
  and AND2_158 (keyinput_Wire_0[26], N146, N483);
  xnor keyGate_0_26(KeyNOTWire_0[11], keyinput26, keyinput_Wire_0[26]);
  not KeyNOTGate_0_11(N512, KeyNOTWire_0[11]);
  and AND2_159 (keyinput_Wire_0[27], N116, N466);
  xnor keyGate_0_27(N513, keyinput27, keyinput_Wire_0[27]);
  and AND2_160 (keyinput_Wire_0[28], N149, N483);
  xor keyGate_0_28(KeyNOTWire_0[12], keyinput28, keyinput_Wire_0[28]);
  not KeyNOTGate_0_12(N514, KeyNOTWire_0[12]);
  and AND2_161 (keyinput_Wire_0[29], N121, N466);
  xor keyGate_0_29(KeyNOTWire_0[13], keyinput29, keyinput_Wire_0[29]);
  not KeyNOTGate_0_13(N515, KeyNOTWire_0[13]);
  and AND2_162 (keyinput_Wire_0[30], N153, N483);
  xnor keyGate_0_30(KeyNOTWire_0[14], keyinput30, keyinput_Wire_0[30]);
  not KeyNOTGate_0_14(N516, KeyNOTWire_0[14]);
  and AND2_163 (keyinput_Wire_0[31], N126, N466);
  xnor keyGate_0_31(KeyNOTWire_0[15], keyinput31, keyinput_Wire_0[31]);
  not KeyNOTGate_0_15(N517, KeyNOTWire_0[15]);
nand NAND2_164 (N518, N130, N492);
or OR2_165 (N519, N130, N492);
nand NAND2_166 (N520, N495, N207);
or OR2_167 (N521, N495, N207);
and AND2_168 (N522, N451, N159);
and AND2_169 (N523, N451, N165);
and AND2_170 (N524, N451, N171);
and AND2_171 (N525, N451, N177);
and AND2_172 (N526, N451, N183);
nand NAND2_173 (N527, N451, N189);
nand NAND2_174 (N528, N451, N195);
nand NAND2_175 (N529, N451, N201);
nand NAND2_176 (N530, N498, N499);
nand NAND2_177 (N533, N500, N501);
nor NOR2_178 (N536, N309, N502);
nor NOR2_179 (N537, N316, N504);
nor NOR2_180 (N538, N317, N506);
nor NOR2_181 (N539, N318, N508);
  nor NOR2_182 (keyinput_Wire_0[32], N510, N511);
  xnor keyGate_0_32(KeyNOTWire_0[16], keyinput32, keyinput_Wire_0[32]);
  not KeyNOTGate_0_16(N540, KeyNOTWire_0[16]);
  nor NOR2_183 (keyinput_Wire_0[33], N512, N513);
  xnor keyGate_0_33(KeyNOTWire_0[17], keyinput33, keyinput_Wire_0[33]);
  not KeyNOTGate_0_17(N541, KeyNOTWire_0[17]);
  nor NOR2_184 (keyinput_Wire_0[34], N514, N515);
  xor keyGate_0_34(KeyNOTWire_0[18], keyinput34, keyinput_Wire_0[34]);
  not KeyNOTGate_0_18(N542, KeyNOTWire_0[18]);
  nor NOR2_185 (keyinput_Wire_0[35], N516, N517);
  xnor keyGate_0_35(KeyNOTWire_0[19], keyinput35, keyinput_Wire_0[35]);
  not KeyNOTGate_0_19(N543, KeyNOTWire_0[19]);
nand NAND2_186 (N544, N518, N519);
nand NAND2_187 (N547, N520, N521);
not NOT1_188 (N550, N530);
not NOT1_189 (N551, N533);
and AND2_190 (N552, N530, N533);
nand NAND2_191 (N553, N536, N503);
nand NAND2_192 (N557, N537, N505);
  nand NAND2_193 (keyinput_Wire_0[36], N538, N507);
  xnor keyGate_0_36(N561, keyinput36, keyinput_Wire_0[36]);
  nand NAND2_194 (keyinput_Wire_0[37], N539, N509);
  xnor keyGate_0_37(KeyNOTWire_0[20], keyinput37, keyinput_Wire_0[37]);
  not KeyNOTGate_0_20(N565, KeyNOTWire_0[20]);
  nand NAND2_195 (keyinput_Wire_0[38], N488, N540);
  xnor keyGate_0_38(N569, keyinput38, keyinput_Wire_0[38]);
  nand NAND2_196 (keyinput_Wire_0[39], N489, N541);
  xor keyGate_0_39(KeyNOTWire_0[21], keyinput39, keyinput_Wire_0[39]);
  not KeyNOTGate_0_21(N573, KeyNOTWire_0[21]);
  nand NAND2_197 (keyinput_Wire_0[40], N490, N542);
  xor keyGate_0_40(KeyNOTWire_0[22], keyinput40, keyinput_Wire_0[40]);
  not KeyNOTGate_0_22(N577, KeyNOTWire_0[22]);
  nand NAND2_198 (keyinput_Wire_0[41], N491, N543);
  xor keyGate_0_41(KeyNOTWire_0[23], keyinput41, keyinput_Wire_0[41]);
  not KeyNOTGate_0_23(N581, KeyNOTWire_0[23]);
not NOT1_199 (N585, N544);
not NOT1_200 (N586, N547);
and AND2_201 (N587, N544, N547);
and AND2_202 (N588, N550, N551);
and AND2_203 (N589, N585, N586);
nand NAND2_204 (N590, N553, N159);
or OR2_205 (N593, N553, N159);
and AND2_206 (N596, N246, N553);
nand NAND2_207 (N597, N557, N165);
or OR2_208 (N600, N557, N165);
and AND2_209 (N605, N246, N557);
nand NAND2_210 (N606, N561, N171);
or OR2_211 (N609, N561, N171);
and AND2_212 (N615, N246, N561);
  nand NAND2_213 (keyinput_Wire_0[42], N565, N177);
  xnor keyGate_0_42(KeyNOTWire_0[24], keyinput42, keyinput_Wire_0[42]);
  not KeyNOTGate_0_24(N616, KeyNOTWire_0[24]);
  or OR2_214 (keyinput_Wire_0[43], N565, N177);
  xnor keyGate_0_43(N619, keyinput43, keyinput_Wire_0[43]);
and AND2_215 (N624, N246, N565);
  nand NAND2_216 (keyinput_Wire_0[44], N569, N183);
  xnor keyGate_0_44(KeyNOTWire_0[25], keyinput44, keyinput_Wire_0[44]);
  not KeyNOTGate_0_25(N625, KeyNOTWire_0[25]);
  or OR2_217 (keyinput_Wire_0[45], N569, N183);
  xnor keyGate_0_45(N628, keyinput45, keyinput_Wire_0[45]);
and AND2_218 (N631, N246, N569);
  nand NAND2_219 (keyinput_Wire_0[46], N573, N189);
  xor keyGate_0_46(KeyNOTWire_0[26], keyinput46, keyinput_Wire_0[46]);
  not KeyNOTGate_0_26(N632, KeyNOTWire_0[26]);
  or OR2_220 (keyinput_Wire_0[47], N573, N189);
  xor keyGate_0_47(N635, keyinput47, keyinput_Wire_0[47]);
and AND2_221 (N640, N246, N573);
  nand NAND2_222 (keyinput_Wire_0[48], N577, N195);
  xnor keyGate_0_48(KeyNOTWire_0[27], keyinput48, keyinput_Wire_0[48]);
  not KeyNOTGate_0_27(N641, KeyNOTWire_0[27]);
  or OR2_223 (keyinput_Wire_0[49], N577, N195);
  xor keyGate_0_49(N644, keyinput49, keyinput_Wire_0[49]);
and AND2_224 (N650, N246, N577);
  nand NAND2_225 (keyinput_Wire_0[50], N581, N201);
  xnor keyGate_0_50(KeyNOTWire_0[28], keyinput50, keyinput_Wire_0[50]);
  not KeyNOTGate_0_28(N651, KeyNOTWire_0[28]);
  or OR2_226 (keyinput_Wire_0[51], N581, N201);
  xnor keyGate_0_51(N654, keyinput51, keyinput_Wire_0[51]);
and AND2_227 (N659, N246, N581);
nor NOR2_228 (N660, N552, N588);
nor NOR2_229 (N661, N587, N589);
not NOT1_230 (N662, N590);
and AND2_231 (N665, N593, N590);
nor NOR2_232 (N669, N596, N522);
not NOT1_233 (N670, N597);
and AND2_234 (N673, N600, N597);
nor NOR2_235 (N677, N605, N523);
not NOT1_236 (N678, N606);
and AND2_237 (N682, N609, N606);
nor NOR2_238 (N686, N615, N524);
not NOT1_239 (N687, N616);
and AND2_240 (N692, N619, N616);
nor NOR2_241 (N696, N624, N525);
  not NOT1_242 (keyinput_Wire_0[52], N625);
  xor keyGate_0_52(KeyNOTWire_0[29], keyinput52, keyinput_Wire_0[52]);
  not KeyNOTGate_0_29(N697, KeyNOTWire_0[29]);
and AND2_243 (N700, N628, N625);
nor NOR2_244 (N704, N631, N526);
  not NOT1_245 (keyinput_Wire_0[53], N632);
  xor keyGate_0_53(KeyNOTWire_0[30], keyinput53, keyinput_Wire_0[53]);
  not KeyNOTGate_0_30(N705, KeyNOTWire_0[30]);
and AND2_246 (N708, N635, N632);
nor NOR2_247 (N712, N337, N640);
  not NOT1_248 (keyinput_Wire_0[54], N641);
  xor keyGate_0_54(N713, keyinput54, keyinput_Wire_0[54]);
and AND2_249 (N717, N644, N641);
nor NOR2_250 (N721, N339, N650);
  not NOT1_251 (keyinput_Wire_0[55], N651);
  xnor keyGate_0_55(KeyNOTWire_0[31], keyinput55, keyinput_Wire_0[55]);
  not KeyNOTGate_0_31(N722, KeyNOTWire_0[31]);
and AND2_252 (N727, N654, N651);
nor NOR2_253 (N731, N341, N659);
nand NAND2_254 (N732, N654, N261);
nand NAND3_255 (N733, N644, N654, N261);
  nand NAND4_256 (keyinput_Wire_0[56], N635, N644, N654, N261);
  xor keyGate_0_56(N734, keyinput56, keyinput_Wire_0[56]);
not NOT1_257 (N735, N662);
and AND2_258 (N736, N228, N665);
and AND2_259 (N737, N237, N662);
not NOT1_260 (N738, N670);
and AND2_261 (N739, N228, N673);
and AND2_262 (N740, N237, N670);
not NOT1_263 (N741, N678);
and AND2_264 (N742, N228, N682);
and AND2_265 (N743, N237, N678);
not NOT1_266 (N744, N687);
and AND2_267 (N745, N228, N692);
and AND2_268 (N746, N237, N687);
  not NOT1_269 (keyinput_Wire_0[57], N697);
  xnor keyGate_0_57(KeyNOTWire_0[32], keyinput57, keyinput_Wire_0[57]);
  not KeyNOTGate_0_32(N747, KeyNOTWire_0[32]);
and AND2_270 (N748, N228, N700);
and AND2_271 (N749, N237, N697);
  not NOT1_272 (keyinput_Wire_0[58], N705);
  xnor keyGate_0_58(KeyNOTWire_0[33], keyinput58, keyinput_Wire_0[58]);
  not KeyNOTGate_0_33(N750, KeyNOTWire_0[33]);
and AND2_273 (N751, N228, N708);
and AND2_274 (N752, N237, N705);
not NOT1_275 (N753, N713);
and AND2_276 (N754, N228, N717);
and AND2_277 (N755, N237, N713);
not NOT1_278 (N756, N722);
nor NOR2_279 (N757, N727, N261);
and AND2_280 (N758, N727, N261);
and AND2_281 (N759, N228, N727);
and AND2_282 (N760, N237, N722);
nand NAND2_283 (N761, N644, N722);
  nand NAND2_284 (keyinput_Wire_0[59], N635, N713);
  xor keyGate_0_59(N762, keyinput59, keyinput_Wire_0[59]);
  nand NAND3_285 (keyinput_Wire_0[60], N635, N644, N722);
  xor keyGate_0_60(KeyNOTWire_0[34], keyinput60, keyinput_Wire_0[60]);
  not KeyNOTGate_0_34(N763, KeyNOTWire_0[34]);
nand NAND2_286 (N764, N609, N687);
nand NAND2_287 (N765, N600, N678);
  nand NAND3_288 (keyinput_Wire_0[61], N600, N609, N687);
  xnor keyGate_0_61(N766, keyinput61, keyinput_Wire_0[61]);
buf BUFF1_289 (N767, N660);
buf BUFF1_290 (N768, N661);
nor NOR2_291 (N769, N736, N737);
nor NOR2_292 (N770, N739, N740);
nor NOR2_293 (N771, N742, N743);
nor NOR2_294 (N772, N745, N746);
  nand NAND4_295 (keyinput_Wire_0[62], N750, N762, N763, N734);
  xor keyGate_0_62(KeyNOTWire_0[35], keyinput62, keyinput_Wire_0[62]);
  not KeyNOTGate_0_35(N773, KeyNOTWire_0[35]);
nor NOR2_296 (N777, N748, N749);
nand NAND3_297 (N778, N753, N761, N733);
nor NOR2_298 (N781, N751, N752);
nand NAND2_299 (N782, N756, N732);
nor NOR2_300 (N785, N754, N755);
nor NOR2_301 (N786, N757, N758);
nor NOR2_302 (N787, N759, N760);
  nor NOR2_303 (keyinput_Wire_0[63], N700, N773);
  xor keyGate_0_63(KeyNOTWire_0[36], keyinput63, keyinput_Wire_0[63]);
  not KeyNOTGate_0_36(N788, KeyNOTWire_0[36]);
  and AND2_304 (keyinput_Wire_0[64], N700, N773);
  xnor keyGate_0_64(N789, keyinput64, keyinput_Wire_0[64]);
  nor NOR2_305 (keyinput_Wire_0[65], N708, N778);
  xnor keyGate_0_65(KeyNOTWire_0[37], keyinput65, keyinput_Wire_0[65]);
  not KeyNOTGate_0_37(N790, KeyNOTWire_0[37]);
  and AND2_306 (keyinput_Wire_0[66], N708, N778);
  xor keyGate_0_66(N791, keyinput66, keyinput_Wire_0[66]);
nor NOR2_307 (N792, N717, N782);
and AND2_308 (N793, N717, N782);
and AND2_309 (N794, N219, N786);
  nand NAND2_310 (keyinput_Wire_0[67], N628, N773);
  xnor keyGate_0_67(KeyNOTWire_0[38], keyinput67, keyinput_Wire_0[67]);
  not KeyNOTGate_0_38(N795, KeyNOTWire_0[38]);
  nand NAND2_311 (keyinput_Wire_0[68], N795, N747);
  xor keyGate_0_68(KeyNOTWire_0[39], keyinput68, keyinput_Wire_0[68]);
  not KeyNOTGate_0_39(N796, KeyNOTWire_0[39]);
  nor NOR2_312 (keyinput_Wire_0[69], N788, N789);
  xor keyGate_0_69(N802, keyinput69, keyinput_Wire_0[69]);
  nor NOR2_313 (keyinput_Wire_0[70], N790, N791);
  xnor keyGate_0_70(KeyNOTWire_0[40], keyinput70, keyinput_Wire_0[70]);
  not KeyNOTGate_0_40(N803, KeyNOTWire_0[40]);
nor NOR2_314 (N804, N792, N793);
nor NOR2_315 (N805, N340, N794);
  nor NOR2_316 (keyinput_Wire_0[71], N692, N796);
  xor keyGate_0_71(N806, keyinput71, keyinput_Wire_0[71]);
  and AND2_317 (keyinput_Wire_0[72], N692, N796);
  xnor keyGate_0_72(KeyNOTWire_0[41], keyinput72, keyinput_Wire_0[72]);
  not KeyNOTGate_0_41(N807, KeyNOTWire_0[41]);
  and AND2_318 (keyinput_Wire_0[73], N219, N802);
  xor keyGate_0_73(N808, keyinput73, keyinput_Wire_0[73]);
  and AND2_319 (keyinput_Wire_0[74], N219, N803);
  xnor keyGate_0_74(KeyNOTWire_0[42], keyinput74, keyinput_Wire_0[74]);
  not KeyNOTGate_0_42(N809, KeyNOTWire_0[42]);
and AND2_320 (N810, N219, N804);
  nand NAND4_321 (keyinput_Wire_0[75], N805, N787, N731, N529);
  xor keyGate_0_75(N811, keyinput75, keyinput_Wire_0[75]);
  nand NAND2_322 (keyinput_Wire_0[76], N619, N796);
  xor keyGate_0_76(N812, keyinput76, keyinput_Wire_0[76]);
  nand NAND3_323 (keyinput_Wire_0[77], N609, N619, N796);
  xnor keyGate_0_77(N813, keyinput77, keyinput_Wire_0[77]);
  nand NAND4_324 (keyinput_Wire_0[78], N600, N609, N619, N796);
  xor keyGate_0_78(N814, keyinput78, keyinput_Wire_0[78]);
  nand NAND4_325 (keyinput_Wire_0[79], N738, N765, N766, N814);
  xor keyGate_0_79(N815, keyinput79, keyinput_Wire_0[79]);
  nand NAND3_326 (keyinput_Wire_0[80], N741, N764, N813);
  xnor keyGate_0_80(KeyNOTWire_0[43], keyinput80, keyinput_Wire_0[80]);
  not KeyNOTGate_0_43(N819, KeyNOTWire_0[43]);
  nand NAND2_327 (keyinput_Wire_0[81], N744, N812);
  xor keyGate_0_81(KeyNOTWire_0[44], keyinput81, keyinput_Wire_0[81]);
  not KeyNOTGate_0_44(N822, KeyNOTWire_0[44]);
  nor NOR2_328 (keyinput_Wire_0[82], N806, N807);
  xor keyGate_0_82(KeyNOTWire_0[45], keyinput82, keyinput_Wire_0[82]);
  not KeyNOTGate_0_45(N825, KeyNOTWire_0[45]);
  nor NOR2_329 (keyinput_Wire_0[83], N335, N808);
  xnor keyGate_0_83(KeyNOTWire_0[46], keyinput83, keyinput_Wire_0[83]);
  not KeyNOTGate_0_46(N826, KeyNOTWire_0[46]);
  nor NOR2_330 (keyinput_Wire_0[84], N336, N809);
  xor keyGate_0_84(N827, keyinput84, keyinput_Wire_0[84]);
nor NOR2_331 (N828, N338, N810);
  not NOT1_332 (keyinput_Wire_0[85], N811);
  xor keyGate_0_85(N829, keyinput85, keyinput_Wire_0[85]);
  nor NOR2_333 (keyinput_Wire_0[86], N665, N815);
  xor keyGate_0_86(KeyNOTWire_0[47], keyinput86, keyinput_Wire_0[86]);
  not KeyNOTGate_0_47(N830, KeyNOTWire_0[47]);
  and AND2_334 (keyinput_Wire_0[87], N665, N815);
  xnor keyGate_0_87(N831, keyinput87, keyinput_Wire_0[87]);
  nor NOR2_335 (keyinput_Wire_0[88], N673, N819);
  xnor keyGate_0_88(N832, keyinput88, keyinput_Wire_0[88]);
  and AND2_336 (keyinput_Wire_0[89], N673, N819);
  xnor keyGate_0_89(N833, keyinput89, keyinput_Wire_0[89]);
  nor NOR2_337 (keyinput_Wire_0[90], N682, N822);
  xor keyGate_0_90(KeyNOTWire_0[48], keyinput90, keyinput_Wire_0[90]);
  not KeyNOTGate_0_48(N834, KeyNOTWire_0[48]);
  and AND2_338 (keyinput_Wire_0[91], N682, N822);
  xnor keyGate_0_91(KeyNOTWire_0[49], keyinput91, keyinput_Wire_0[91]);
  not KeyNOTGate_0_49(N835, KeyNOTWire_0[49]);
  and AND2_339 (keyinput_Wire_0[92], N219, N825);
  xnor keyGate_0_92(KeyNOTWire_0[50], keyinput92, keyinput_Wire_0[92]);
  not KeyNOTGate_0_50(N836, KeyNOTWire_0[50]);
  nand NAND3_340 (keyinput_Wire_0[93], N826, N777, N704);
  xor keyGate_0_93(N837, keyinput93, keyinput_Wire_0[93]);
  nand NAND4_341 (keyinput_Wire_0[94], N827, N781, N712, N527);
  xnor keyGate_0_94(N838, keyinput94, keyinput_Wire_0[94]);
  nand NAND4_342 (keyinput_Wire_0[95], N828, N785, N721, N528);
  xnor keyGate_0_95(N839, keyinput95, keyinput_Wire_0[95]);
  not NOT1_343 (keyinput_Wire_0[96], N829);
  xnor keyGate_0_96(KeyNOTWire_0[51], keyinput96, keyinput_Wire_0[96]);
  not KeyNOTGate_0_51(N840, KeyNOTWire_0[51]);
  nand NAND2_344 (keyinput_Wire_0[97], N815, N593);
  xnor keyGate_0_97(KeyNOTWire_0[52], keyinput97, keyinput_Wire_0[97]);
  not KeyNOTGate_0_52(N841, KeyNOTWire_0[52]);
  nor NOR2_345 (keyinput_Wire_0[98], N830, N831);
  xor keyGate_0_98(N842, keyinput98, keyinput_Wire_0[98]);
  nor NOR2_346 (keyinput_Wire_0[99], N832, N833);
  xnor keyGate_0_99(N843, keyinput99, keyinput_Wire_0[99]);
  nor NOR2_347 (keyinput_Wire_0[100], N834, N835);
  xor keyGate_0_100(N844, keyinput100, keyinput_Wire_0[100]);
  nor NOR2_348 (keyinput_Wire_0[101], N334, N836);
  xor keyGate_0_101(KeyNOTWire_0[53], keyinput101, keyinput_Wire_0[101]);
  not KeyNOTGate_0_53(N845, KeyNOTWire_0[53]);
  not NOT1_349 (keyinput_Wire_0[102], N837);
  xnor keyGate_0_102(KeyNOTWire_0[54], keyinput102, keyinput_Wire_0[102]);
  not KeyNOTGate_0_54(N846, KeyNOTWire_0[54]);
  not NOT1_350 (keyinput_Wire_0[103], N838);
  xnor keyGate_0_103(KeyNOTWire_0[55], keyinput103, keyinput_Wire_0[103]);
  not KeyNOTGate_0_55(N847, KeyNOTWire_0[55]);
  not NOT1_351 (keyinput_Wire_0[104], N839);
  xnor keyGate_0_104(N848, keyinput104, keyinput_Wire_0[104]);
  and AND2_352 (keyinput_Wire_0[105], N735, N841);
  xnor keyGate_0_105(N849, keyinput105, keyinput_Wire_0[105]);
buf BUFF1_353 (N850, N840);
  and AND2_354 (keyinput_Wire_0[106], N219, N842);
  xor keyGate_0_106(KeyNOTWire_0[56], keyinput106, keyinput_Wire_0[106]);
  not KeyNOTGate_0_56(N851, KeyNOTWire_0[56]);
  and AND2_355 (keyinput_Wire_0[107], N219, N843);
  xnor keyGate_0_107(KeyNOTWire_0[57], keyinput107, keyinput_Wire_0[107]);
  not KeyNOTGate_0_57(N852, KeyNOTWire_0[57]);
  and AND2_356 (keyinput_Wire_0[108], N219, N844);
  xor keyGate_0_108(KeyNOTWire_0[58], keyinput108, keyinput_Wire_0[108]);
  not KeyNOTGate_0_58(N853, KeyNOTWire_0[58]);
  nand NAND3_357 (keyinput_Wire_0[109], N845, N772, N696);
  xnor keyGate_0_109(KeyNOTWire_0[59], keyinput109, keyinput_Wire_0[109]);
  not KeyNOTGate_0_59(N854, KeyNOTWire_0[59]);
  not NOT1_358 (keyinput_Wire_0[110], N846);
  xnor keyGate_0_110(KeyNOTWire_0[60], keyinput110, keyinput_Wire_0[110]);
  not KeyNOTGate_0_60(N855, KeyNOTWire_0[60]);
  not NOT1_359 (keyinput_Wire_0[111], N847);
  xnor keyGate_0_111(N856, keyinput111, keyinput_Wire_0[111]);
  not NOT1_360 (keyinput_Wire_0[112], N848);
  xor keyGate_0_112(KeyNOTWire_0[61], keyinput112, keyinput_Wire_0[112]);
  not KeyNOTGate_0_61(N857, KeyNOTWire_0[61]);
  not NOT1_361 (keyinput_Wire_0[113], N849);
  xnor keyGate_0_113(N858, keyinput113, keyinput_Wire_0[113]);
  nor NOR2_362 (keyinput_Wire_0[114], N417, N851);
  xor keyGate_0_114(N859, keyinput114, keyinput_Wire_0[114]);
  nor NOR2_363 (keyinput_Wire_0[115], N332, N852);
  xor keyGate_0_115(N860, keyinput115, keyinput_Wire_0[115]);
  nor NOR2_364 (keyinput_Wire_0[116], N333, N853);
  xnor keyGate_0_116(KeyNOTWire_0[62], keyinput116, keyinput_Wire_0[116]);
  not KeyNOTGate_0_62(N861, KeyNOTWire_0[62]);
  not NOT1_365 (keyinput_Wire_0[117], N854);
  xnor keyGate_0_117(N862, keyinput117, keyinput_Wire_0[117]);
buf BUFF1_366 (N863, N855);
buf BUFF1_367 (N864, N856);
buf BUFF1_368 (N865, N857);
  buf BUFF1_369 (keyinput_Wire_1, N858);
  xor keyGate_1_9(N866, KeyWire_0_2, keyinput_Wire_1);
  nand NAND3_370 (keyinput_Wire_0[118], N859, N769, N669);
  xor keyGate_0_118(KeyNOTWire_0[63], keyinput118, keyinput_Wire_0[118]);
  not KeyNOTGate_0_63(N867, KeyNOTWire_0[63]);
  nand NAND3_371 (keyinput_Wire_0[119], N860, N770, N677);
  xor keyGate_0_119(KeyNOTWire_0[64], keyinput119, keyinput_Wire_0[119]);
  not KeyNOTGate_0_64(N868, KeyNOTWire_0[64]);
  nand NAND3_372 (keyinput_Wire_0[120], N861, N771, N686);
  xor keyGate_0_120(N869, keyinput120, keyinput_Wire_0[120]);
  not NOT1_373 (keyinput_Wire_0[121], N862);
  xor keyGate_0_121(KeyNOTWire_0[65], keyinput121, keyinput_Wire_0[121]);
  not KeyNOTGate_0_65(N870, KeyNOTWire_0[65]);
  not NOT1_374 (keyinput_Wire_0[122], N867);
  xnor keyGate_0_122(KeyNOTWire_0[66], keyinput122, keyinput_Wire_0[122]);
  not KeyNOTGate_0_66(N871, KeyNOTWire_0[66]);
  not NOT1_375 (keyinput_Wire_0[123], N868);
  xor keyGate_0_123(N872, keyinput123, keyinput_Wire_0[123]);
  not NOT1_376 (keyinput_Wire_0[124], N869);
  xor keyGate_0_124(N873, keyinput124, keyinput_Wire_0[124]);
buf BUFF1_377 (N874, N870);
  not NOT1_378 (keyinput_Wire_0[125], N871);
  xor keyGate_0_125(N875, keyinput125, keyinput_Wire_0[125]);
  not NOT1_379 (keyinput_Wire_0[126], N872);
  xor keyGate_0_126(N876, keyinput126, keyinput_Wire_0[126]);
  not NOT1_380 (keyinput_Wire_0[127], N873);
  xnor keyGate_0_127(N877, keyinput127, keyinput_Wire_0[127]);
buf BUFF1_381 (KeyWire_0_1, N875);
  xor flip_it (N878, KeyWire_0_1, KeyWire_0_2 );
buf BUFF1_382 (N879, N876);
buf BUFF1_383 (N880, N877);

AntiSAT some_name( KeyWire_0_2, N86, N17, N42, N156, N237, N260, N255, N177, N87, N171, N126, N36, N88, N143, N165, N29, N90, N26, N183, N246, N116, N89, N152, N72, N80, N189, N219, N267, N195, N59, N51, N111, N207, N159, N228, N68, N96, N13, N130, N149, N75, N210, N85, N201, N91, N259, N73, N74, N106, N153, N138, N55, N101, N268, N1, N121, N146, N8, N261, N135, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, keyinput245, keyinput246, keyinput247,
       keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
       keyinput253, keyinput254, keyinput255, keyinput256, keyinput257,
       keyinput258, keyinput259, keyinput260, keyinput261, keyinput262,
       keyinput263, keyinput264, keyinput265, keyinput266, keyinput267,
       keyinput268, keyinput269, keyinput270, keyinput271, keyinput272,
       keyinput273, keyinput274, keyinput275, keyinput276, keyinput277,
       keyinput278, keyinput279, keyinput280, keyinput281, keyinput282,
       keyinput283, keyinput284, keyinput285, keyinput286, keyinput287,
       keyinput288, keyinput289, keyinput290, keyinput291, keyinput292,
       keyinput293, keyinput294, keyinput295, keyinput296, keyinput297,
       keyinput298, keyinput299, keyinput300, keyinput301, keyinput302,
       keyinput303, keyinput304, keyinput305, keyinput306, keyinput307);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N86, N17, N42, N156, N237, N260, N255, N177, N87, N171, N126, N36, N88, N143, N165, N29, N90, N26, N183, N246, N116, N89, N152, N72, N80, N189, N219, N267, N195, N59, N51, N111, N207, N159, N228, N68, N96, N13, N130, N149, N75, N210, N85, N201, N91, N259, N73, N74, N106, N153, N138, N55, N101, N268, N1, N121, N146, N8, N261, N135, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, keyinput245, keyinput246, keyinput247 ,
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
        keyinput253, keyinput254, keyinput255, keyinput256, keyinput257,
        keyinput258, keyinput259, keyinput260, keyinput261, keyinput262,
        keyinput263, keyinput264, keyinput265, keyinput266, keyinput267,
        keyinput268, keyinput269, keyinput270, keyinput271, keyinput272,
        keyinput273, keyinput274, keyinput275, keyinput276, keyinput277,
        keyinput278, keyinput279, keyinput280, keyinput281, keyinput282,
        keyinput283, keyinput284, keyinput285, keyinput286, keyinput287,
        keyinput288, keyinput289, keyinput290, keyinput291, keyinput292,
        keyinput293, keyinput294, keyinput295, keyinput296, keyinput297,
        keyinput298, keyinput299, keyinput300, keyinput301, keyinput302,
        keyinput303, keyinput304, keyinput305, keyinput306, keyinput307);

  input keyinput248, keyinput249, keyinput250, keyinput251, keyinput252;
  input keyinput253, keyinput254, keyinput255, keyinput256, keyinput257;
  input keyinput258, keyinput259, keyinput260, keyinput261, keyinput262;
  input keyinput263, keyinput264, keyinput265, keyinput266, keyinput267;
  input keyinput268, keyinput269, keyinput270, keyinput271, keyinput272;
  input keyinput273, keyinput274, keyinput275, keyinput276, keyinput277;
  input keyinput278, keyinput279, keyinput280, keyinput281, keyinput282;
  input keyinput283, keyinput284, keyinput285, keyinput286, keyinput287;
  input keyinput288, keyinput289, keyinput290, keyinput291, keyinput292;
  input keyinput293, keyinput294, keyinput295, keyinput296, keyinput297;
  input keyinput298, keyinput299, keyinput300, keyinput301, keyinput302;
  input keyinput303, keyinput304, keyinput305, keyinput306, keyinput307;

  wire [0:59] keyNTin_Wire_1;
  wire [0:30] KeyNOTWire_1;

  input N86, N17, N42, N156, N237, N260, N255, N177, N87, N171, N126, N36, N88, N143, N165, N29, N90, N26, N183, N246, N116, N89, N152, N72, N80, N189, N219, N267, N195, N59, N51, N111, N207, N159, N228, N68, N96, N13, N130, N149, N75, N210, N85, N201, N91, N259, N73, N74, N106, N153, N138, N55, N101, N268, N1, N121, N146, N8, N261, N135;
  input keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, keyinput245, keyinput246, keyinput247;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83, newWire_84, newWire_85, newWire_86, newWire_87, newWire_88, newWire_89, newWire_90, newWire_91, newWire_92, newWire_93, newWire_94, newWire_95, newWire_96, newWire_97, newWire_98, newWire_99, newWire_100, newWire_101, newWire_102, newWire_103, newWire_104, newWire_105, newWire_106, newWire_107, newWire_108, newWire_109, newWire_110, newWire_111, newWire_112, newWire_113, newWire_114, newWire_115, newWire_116, newWire_117, newWire_118, newWire_119, newWire_120, newWire_121 ;

  xnor KeyGate0 (keyNTin_Wire_1[0], N86, keyinput128);
  xor keyNTinGate_1_0(newWire_0, keyinput248, keyNTin_Wire_1[0]);
  xnor KeyGate1 (newWire_1, N17, keyinput129);
  xnor KeyGate2 (keyNTin_Wire_1[1], N42, keyinput130);
  xnor keyNTinGate_1_1(newWire_2, keyinput249, keyNTin_Wire_1[1]);
  xnor KeyGate3 (newWire_3, N156, keyinput131);
  xnor KeyGate4 (newWire_4, N237, keyinput132);
  xor  KeyGate5 (newWire_5, N260, keyinput133);
  xnor KeyGate6 (keyNTin_Wire_1[2], N255, keyinput134);
  xnor keyNTinGate_1_2(newWire_6, keyinput250, keyNTin_Wire_1[2]);
  xnor KeyGate7 (newWire_7, N177, keyinput135);
  xnor KeyGate8 (keyNTin_Wire_1[3], N87, keyinput136);
  xnor keyNTinGate_1_3(newWire_8, keyinput251, keyNTin_Wire_1[3]);
  xor  KeyGate9 (newWire_9, N171, keyinput137);
  xor  KeyGate10 (keyNTin_Wire_1[4], N126, keyinput138);
  xnor keyNTinGate_1_4(KeyNOTWire_1[0], keyinput252, keyNTin_Wire_1[4]);
  not KeyNOTGate_1_0(newWire_10, KeyNOTWire_1[0]);
  xor  KeyGate11 (keyNTin_Wire_1[5], N36, keyinput139);
  xnor keyNTinGate_1_5(KeyNOTWire_1[1], keyinput253, keyNTin_Wire_1[5]);
  not KeyNOTGate_1_1(newWire_11, KeyNOTWire_1[1]);
  xor  KeyGate12 (newWire_12, N88, keyinput140);
  xnor KeyGate13 (keyNTin_Wire_1[6], N143, keyinput141);
  xnor keyNTinGate_1_6(KeyNOTWire_1[2], keyinput254, keyNTin_Wire_1[6]);
  not KeyNOTGate_1_2(newWire_13, KeyNOTWire_1[2]);
  xnor KeyGate14 (keyNTin_Wire_1[7], N165, keyinput142);
  xnor keyNTinGate_1_7(newWire_14, keyinput255, keyNTin_Wire_1[7]);
  xnor KeyGate15 (newWire_15, N29, keyinput143);
  xor  KeyGate16 (keyNTin_Wire_1[8], N90, keyinput144);
  xnor keyNTinGate_1_8(KeyNOTWire_1[3], keyinput256, keyNTin_Wire_1[8]);
  not KeyNOTGate_1_3(newWire_16, KeyNOTWire_1[3]);
  xnor KeyGate17 (keyNTin_Wire_1[9], N26, keyinput145);
  xor keyNTinGate_1_9(newWire_17, keyinput257, keyNTin_Wire_1[9]);
  xnor KeyGate18 (newWire_18, N183, keyinput146);
  xnor KeyGate19 (keyNTin_Wire_1[10], N246, keyinput147);
  xnor keyNTinGate_1_10(KeyNOTWire_1[4], keyinput258, keyNTin_Wire_1[10]);
  not KeyNOTGate_1_4(newWire_19, KeyNOTWire_1[4]);
  xnor KeyGate20 (newWire_20, N116, keyinput148);
  xnor KeyGate21 (keyNTin_Wire_1[11], N89, keyinput149);
  xor keyNTinGate_1_11(KeyNOTWire_1[5], keyinput259, keyNTin_Wire_1[11]);
  not KeyNOTGate_1_5(newWire_21, KeyNOTWire_1[5]);
  xor  KeyGate22 (newWire_22, N152, keyinput150);
  xnor KeyGate23 (keyNTin_Wire_1[12], N72, keyinput151);
  xnor keyNTinGate_1_12(KeyNOTWire_1[6], keyinput260, keyNTin_Wire_1[12]);
  not KeyNOTGate_1_6(newWire_23, KeyNOTWire_1[6]);
  xnor KeyGate24 (keyNTin_Wire_1[13], N80, keyinput152);
  xor keyNTinGate_1_13(newWire_24, keyinput261, keyNTin_Wire_1[13]);
  xnor KeyGate25 (newWire_25, N189, keyinput153);
  xor  KeyGate26 (newWire_26, N219, keyinput154);
  xor  KeyGate27 (keyNTin_Wire_1[14], N267, keyinput155);
  xor keyNTinGate_1_14(newWire_27, keyinput262, keyNTin_Wire_1[14]);
  xnor KeyGate28 (keyNTin_Wire_1[15], N195, keyinput156);
  xor keyNTinGate_1_15(KeyNOTWire_1[7], keyinput263, keyNTin_Wire_1[15]);
  not KeyNOTGate_1_7(newWire_28, KeyNOTWire_1[7]);
  xnor KeyGate29 (keyNTin_Wire_1[16], N59, keyinput157);
  xor keyNTinGate_1_16(KeyNOTWire_1[8], keyinput264, keyNTin_Wire_1[16]);
  not KeyNOTGate_1_8(newWire_29, KeyNOTWire_1[8]);
  xor  KeyGate30 (newWire_30, N51, keyinput158);
  xor  KeyGate31 (newWire_31, N111, keyinput159);
  xnor KeyGate32 (newWire_32, N207, keyinput160);
  xnor KeyGate33 (newWire_33, N159, keyinput161);
  xnor KeyGate34 (keyNTin_Wire_1[17], N228, keyinput162);
  xnor keyNTinGate_1_17(newWire_34, keyinput265, keyNTin_Wire_1[17]);
  xnor KeyGate35 (newWire_35, N68, keyinput163);
  xnor KeyGate36 (keyNTin_Wire_1[18], N96, keyinput164);
  xor keyNTinGate_1_18(newWire_36, keyinput266, keyNTin_Wire_1[18]);
  xnor KeyGate37 (keyNTin_Wire_1[19], N13, keyinput165);
  xnor keyNTinGate_1_19(KeyNOTWire_1[9], keyinput267, keyNTin_Wire_1[19]);
  not KeyNOTGate_1_9(newWire_37, KeyNOTWire_1[9]);
  xnor KeyGate38 (keyNTin_Wire_1[20], N130, keyinput166);
  xnor keyNTinGate_1_20(KeyNOTWire_1[10], keyinput268, keyNTin_Wire_1[20]);
  not KeyNOTGate_1_10(newWire_38, KeyNOTWire_1[10]);
  xor  KeyGate39 (keyNTin_Wire_1[21], N149, keyinput167);
  xor keyNTinGate_1_21(newWire_39, keyinput269, keyNTin_Wire_1[21]);
  xor  KeyGate40 (keyNTin_Wire_1[22], N75, keyinput168);
  xor keyNTinGate_1_22(KeyNOTWire_1[11], keyinput270, keyNTin_Wire_1[22]);
  not KeyNOTGate_1_11(newWire_40, KeyNOTWire_1[11]);
  xnor KeyGate41 (keyNTin_Wire_1[23], N210, keyinput169);
  xnor keyNTinGate_1_23(KeyNOTWire_1[12], keyinput271, keyNTin_Wire_1[23]);
  not KeyNOTGate_1_12(newWire_41, KeyNOTWire_1[12]);
  xnor KeyGate42 (keyNTin_Wire_1[24], N85, keyinput170);
  xnor keyNTinGate_1_24(newWire_42, keyinput272, keyNTin_Wire_1[24]);
  xnor KeyGate43 (keyNTin_Wire_1[25], N201, keyinput171);
  xor keyNTinGate_1_25(KeyNOTWire_1[13], keyinput273, keyNTin_Wire_1[25]);
  not KeyNOTGate_1_13(newWire_43, KeyNOTWire_1[13]);
  xnor KeyGate44 (newWire_44, N91, keyinput172);
  xor  KeyGate45 (keyNTin_Wire_1[26], N259, keyinput173);
  xor keyNTinGate_1_26(newWire_45, keyinput274, keyNTin_Wire_1[26]);
  xor  KeyGate46 (keyNTin_Wire_1[27], N73, keyinput174);
  xnor keyNTinGate_1_27(KeyNOTWire_1[14], keyinput275, keyNTin_Wire_1[27]);
  not KeyNOTGate_1_14(newWire_46, KeyNOTWire_1[14]);
  xnor KeyGate47 (keyNTin_Wire_1[28], N74, keyinput175);
  xor keyNTinGate_1_28(KeyNOTWire_1[15], keyinput276, keyNTin_Wire_1[28]);
  not KeyNOTGate_1_15(newWire_47, KeyNOTWire_1[15]);
  xor  KeyGate48 (keyNTin_Wire_1[29], N106, keyinput176);
  xnor keyNTinGate_1_29(KeyNOTWire_1[16], keyinput277, keyNTin_Wire_1[29]);
  not KeyNOTGate_1_16(newWire_48, KeyNOTWire_1[16]);
  xnor KeyGate49 (newWire_49, N153, keyinput177);
  xnor KeyGate50 (keyNTin_Wire_1[30], N138, keyinput178);
  xor keyNTinGate_1_30(newWire_50, keyinput278, keyNTin_Wire_1[30]);
  xor  KeyGate51 (newWire_51, N55, keyinput179);
  xor  KeyGate52 (keyNTin_Wire_1[31], N101, keyinput180);
  xnor keyNTinGate_1_31(newWire_52, keyinput279, keyNTin_Wire_1[31]);
  xnor KeyGate53 (newWire_53, N268, keyinput181);
  xnor KeyGate54 (newWire_54, N1, keyinput182);
  xnor KeyGate55 (newWire_55, N121, keyinput183);
  xor  KeyGate56 (newWire_56, N146, keyinput184);
  xnor KeyGate57 (keyNTin_Wire_1[32], N8, keyinput185);
  xnor keyNTinGate_1_32(KeyNOTWire_1[17], keyinput280, keyNTin_Wire_1[32]);
  not KeyNOTGate_1_17(newWire_57, KeyNOTWire_1[17]);
  xnor KeyGate58 (newWire_58, N261, keyinput186);
  xnor KeyGate59 (newWire_59, N135, keyinput187);
  xor  KeyGate60 (keyNTin_Wire_1[33], N86, keyinput188);
  xnor keyNTinGate_1_33(newWire_60, keyinput281, keyNTin_Wire_1[33]);
  xnor KeyGate61 (keyNTin_Wire_1[34], N17, keyinput189);
  xor keyNTinGate_1_34(newWire_61, keyinput282, keyNTin_Wire_1[34]);
  xor  KeyGate62 (newWire_62, N42, keyinput190);
  xor  KeyGate63 (keyNTin_Wire_1[35], N156, keyinput191);
  xnor keyNTinGate_1_35(KeyNOTWire_1[18], keyinput283, keyNTin_Wire_1[35]);
  not KeyNOTGate_1_18(newWire_63, KeyNOTWire_1[18]);
  xor  KeyGate64 (keyNTin_Wire_1[36], N237, keyinput192);
  xor keyNTinGate_1_36(newWire_64, keyinput284, keyNTin_Wire_1[36]);
  xnor KeyGate65 (newWire_65, N260, keyinput193);
  xnor KeyGate66 (newWire_66, N255, keyinput194);
  xnor KeyGate67 (newWire_67, N177, keyinput195);
  xor  KeyGate68 (keyNTin_Wire_1[37], N87, keyinput196);
  xor keyNTinGate_1_37(newWire_68, keyinput285, keyNTin_Wire_1[37]);
  xor  KeyGate69 (newWire_69, N171, keyinput197);
  xnor KeyGate70 (newWire_70, N126, keyinput198);
  xnor KeyGate71 (newWire_71, N36, keyinput199);
  xor  KeyGate72 (newWire_72, N88, keyinput200);
  xnor KeyGate73 (newWire_73, N143, keyinput201);
  xnor KeyGate74 (keyNTin_Wire_1[38], N165, keyinput202);
  xnor keyNTinGate_1_38(newWire_74, keyinput286, keyNTin_Wire_1[38]);
  xnor KeyGate75 (keyNTin_Wire_1[39], N29, keyinput203);
  xor keyNTinGate_1_39(KeyNOTWire_1[19], keyinput287, keyNTin_Wire_1[39]);
  not KeyNOTGate_1_19(newWire_75, KeyNOTWire_1[19]);
  xor  KeyGate76 (keyNTin_Wire_1[40], N90, keyinput204);
  xor keyNTinGate_1_40(KeyNOTWire_1[20], keyinput288, keyNTin_Wire_1[40]);
  not KeyNOTGate_1_20(newWire_76, KeyNOTWire_1[20]);
  xor  KeyGate77 (newWire_77, N26, keyinput205);
  xnor KeyGate78 (newWire_78, N183, keyinput206);
  xnor KeyGate79 (newWire_79, N246, keyinput207);
  xor  KeyGate80 (newWire_80, N116, keyinput208);
  xnor KeyGate81 (keyNTin_Wire_1[41], N89, keyinput209);
  xnor keyNTinGate_1_41(KeyNOTWire_1[21], keyinput289, keyNTin_Wire_1[41]);
  not KeyNOTGate_1_21(newWire_81, KeyNOTWire_1[21]);
  xor  KeyGate82 (keyNTin_Wire_1[42], N152, keyinput210);
  xor keyNTinGate_1_42(KeyNOTWire_1[22], keyinput290, keyNTin_Wire_1[42]);
  not KeyNOTGate_1_22(newWire_82, KeyNOTWire_1[22]);
  xnor KeyGate83 (keyNTin_Wire_1[43], N72, keyinput211);
  xor keyNTinGate_1_43(newWire_83, keyinput291, keyNTin_Wire_1[43]);
  xnor KeyGate84 (newWire_84, N80, keyinput212);
  xor  KeyGate85 (newWire_85, N189, keyinput213);
  xnor KeyGate86 (newWire_86, N219, keyinput214);
  xor  KeyGate87 (keyNTin_Wire_1[44], N267, keyinput215);
  xnor keyNTinGate_1_44(newWire_87, keyinput292, keyNTin_Wire_1[44]);
  xnor KeyGate88 (newWire_88, N195, keyinput216);
  xnor KeyGate89 (keyNTin_Wire_1[45], N59, keyinput217);
  xnor keyNTinGate_1_45(newWire_89, keyinput293, keyNTin_Wire_1[45]);
  xor  KeyGate90 (keyNTin_Wire_1[46], N51, keyinput218);
  xor keyNTinGate_1_46(newWire_90, keyinput294, keyNTin_Wire_1[46]);
  xnor KeyGate91 (keyNTin_Wire_1[47], N111, keyinput219);
  xnor keyNTinGate_1_47(KeyNOTWire_1[23], keyinput295, keyNTin_Wire_1[47]);
  not KeyNOTGate_1_23(newWire_91, KeyNOTWire_1[23]);
  xnor KeyGate92 (newWire_92, N207, keyinput220);
  xnor KeyGate93 (newWire_93, N159, keyinput221);
  xor  KeyGate94 (newWire_94, N228, keyinput222);
  xnor KeyGate95 (keyNTin_Wire_1[48], N68, keyinput223);
  xnor keyNTinGate_1_48(newWire_95, keyinput296, keyNTin_Wire_1[48]);
  xor  KeyGate96 (keyNTin_Wire_1[49], N96, keyinput224);
  xor keyNTinGate_1_49(newWire_96, keyinput297, keyNTin_Wire_1[49]);
  xnor KeyGate97 (newWire_97, N13, keyinput225);
  xnor KeyGate98 (newWire_98, N130, keyinput226);
  xnor KeyGate99 (newWire_99, N149, keyinput227);
  xor  KeyGate100 (keyNTin_Wire_1[50], N75, keyinput228);
  xnor keyNTinGate_1_50(KeyNOTWire_1[24], keyinput298, keyNTin_Wire_1[50]);
  not KeyNOTGate_1_24(newWire_100, KeyNOTWire_1[24]);
  xor  KeyGate101 (keyNTin_Wire_1[51], N210, keyinput229);
  xor keyNTinGate_1_51(newWire_101, keyinput299, keyNTin_Wire_1[51]);
  xor  KeyGate102 (keyNTin_Wire_1[52], N85, keyinput230);
  xor keyNTinGate_1_52(newWire_102, keyinput300, keyNTin_Wire_1[52]);
  xnor KeyGate103 (keyNTin_Wire_1[53], N201, keyinput231);
  xnor keyNTinGate_1_53(KeyNOTWire_1[25], keyinput301, keyNTin_Wire_1[53]);
  not KeyNOTGate_1_25(newWire_103, KeyNOTWire_1[25]);
  xor  KeyGate104 (newWire_104, N91, keyinput232);
  xor  KeyGate105 (newWire_105, N259, keyinput233);
  xnor KeyGate106 (newWire_106, N73, keyinput234);
  xor  KeyGate107 (newWire_107, N74, keyinput235);
  xnor KeyGate108 (newWire_108, N106, keyinput236);
  xnor KeyGate109 (keyNTin_Wire_1[54], N153, keyinput237);
  xnor keyNTinGate_1_54(KeyNOTWire_1[26], keyinput302, keyNTin_Wire_1[54]);
  not KeyNOTGate_1_26(newWire_109, KeyNOTWire_1[26]);
  xor  KeyGate110 (newWire_110, N138, keyinput238);
  xnor KeyGate111 (newWire_111, N55, keyinput239);
  xor  KeyGate112 (keyNTin_Wire_1[55], N101, keyinput240);
  xnor keyNTinGate_1_55(newWire_112, keyinput303, keyNTin_Wire_1[55]);
  xor  KeyGate113 (keyNTin_Wire_1[56], N268, keyinput241);
  xnor keyNTinGate_1_56(KeyNOTWire_1[27], keyinput304, keyNTin_Wire_1[56]);
  not KeyNOTGate_1_27(newWire_113, KeyNOTWire_1[27]);
  xor  KeyGate114 (newWire_114, N1, keyinput242);
  xor  KeyGate115 (newWire_115, N121, keyinput243);
  xor  KeyGate116 (newWire_116, N146, keyinput244);
  xnor KeyGate117 (keyNTin_Wire_1[57], N8, keyinput245);
  xnor keyNTinGate_1_57(KeyNOTWire_1[28], keyinput305, keyNTin_Wire_1[57]);
  not KeyNOTGate_1_28(newWire_117, KeyNOTWire_1[28]);
  xor  KeyGate118 (keyNTin_Wire_1[58], N261, keyinput246);
  xnor keyNTinGate_1_58(KeyNOTWire_1[29], keyinput306, keyNTin_Wire_1[58]);
  not KeyNOTGate_1_29(newWire_118, KeyNOTWire_1[29]);
  xor  KeyGate119 (keyNTin_Wire_1[59], N135, keyinput247);
  xor keyNTinGate_1_59(KeyNOTWire_1[30], keyinput307, keyNTin_Wire_1[59]);
  not KeyNOTGate_1_30(newWire_119, KeyNOTWire_1[30]);
  and some_function (newWire_120, newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59 );
  nand compl_function (newWire_121, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83, newWire_84, newWire_85, newWire_86, newWire_87, newWire_88, newWire_89, newWire_90, newWire_91, newWire_92, newWire_93, newWire_94, newWire_95, newWire_96, newWire_97, newWire_98, newWire_99, newWire_100, newWire_101, newWire_102, newWire_103, newWire_104, newWire_105, newWire_106, newWire_107, newWire_108, newWire_109, newWire_110, newWire_111, newWire_112, newWire_113, newWire_114, newWire_115, newWire_116, newWire_117, newWire_118, newWire_119);
  and finalAND (KeyWire_0_2, newWire_120, newWire_121);

endmodule /* AntiSAT */
