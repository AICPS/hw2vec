`timescale 1ns / 1ps
// Verilog
// c880
// Ninputs 60
// Noutputs 26
// NtotalGates 383
// NAND4 13
// AND3 12
// NAND2 60
// NAND3 14
// AND2 105
// OR2 29
// NOT1 63
// NOR2 61
// BUFF1 26

module top (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
                  N865,N866,N874,N878,N879,N880,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
        keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
                  keyinput125, keyinput126, keyinput127,
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202,
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207,
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212,
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217,
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222,
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227,
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232,
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237,
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242,
                  keyinput243, keyinput244, keyinput245, keyinput246, keyinput247,
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
        keyinput253, keyinput254, keyinput255, keyinput256, keyinput257,
        keyinput258, keyinput259, keyinput260, keyinput261, keyinput262,
        keyinput263, keyinput264, keyinput265, keyinput266, keyinput267,
        keyinput268, keyinput269, keyinput270, keyinput271, keyinput272,
        keyinput273, keyinput274, keyinput275, keyinput276, keyinput277,
        keyinput278, keyinput279, keyinput280, keyinput281, keyinput282,
        keyinput283, keyinput284, keyinput285, keyinput286, keyinput287,
        keyinput288, keyinput289, keyinput290, keyinput291, keyinput292,
        keyinput293, keyinput294, keyinput295, keyinput296, keyinput297,
        keyinput298, keyinput299, keyinput300, keyinput301, keyinput302,
        keyinput303, keyinput304, keyinput305, keyinput306, keyinput307);

  input keyinput248, keyinput249, keyinput250, keyinput251, keyinput252;
  input keyinput253, keyinput254, keyinput255, keyinput256, keyinput257;
  input keyinput258, keyinput259, keyinput260, keyinput261, keyinput262;
  input keyinput263, keyinput264, keyinput265, keyinput266, keyinput267;
  input keyinput268, keyinput269, keyinput270, keyinput271, keyinput272;
  input keyinput273, keyinput274, keyinput275, keyinput276, keyinput277;
  input keyinput278, keyinput279, keyinput280, keyinput281, keyinput282;
  input keyinput283, keyinput284, keyinput285, keyinput286, keyinput287;
  input keyinput288, keyinput289, keyinput290, keyinput291, keyinput292;
  input keyinput293, keyinput294, keyinput295, keyinput296, keyinput297;
  input keyinput298, keyinput299, keyinput300, keyinput301, keyinput302;
  input keyinput303, keyinput304, keyinput305, keyinput306, keyinput307;


  input keyinput128, keyinput129, keyinput130, keyinput131, keyinput132;
  input keyinput133, keyinput134, keyinput135, keyinput136, keyinput137;
  input keyinput138, keyinput139, keyinput140, keyinput141, keyinput142;
  input keyinput143, keyinput144, keyinput145, keyinput146, keyinput147;
  input keyinput148, keyinput149, keyinput150, keyinput151, keyinput152;
  input keyinput153, keyinput154, keyinput155, keyinput156, keyinput157;
  input keyinput158, keyinput159, keyinput160, keyinput161, keyinput162;
  input keyinput163, keyinput164, keyinput165, keyinput166, keyinput167;
  input keyinput168, keyinput169, keyinput170, keyinput171, keyinput172;
  input keyinput173, keyinput174, keyinput175, keyinput176, keyinput177;
  input keyinput178, keyinput179, keyinput180, keyinput181, keyinput182;
  input keyinput183, keyinput184, keyinput185, keyinput186, keyinput187;
  input keyinput188, keyinput189, keyinput190, keyinput191, keyinput192;
  input keyinput193, keyinput194, keyinput195, keyinput196, keyinput197;
  input keyinput198, keyinput199, keyinput200, keyinput201, keyinput202;
  input keyinput203, keyinput204, keyinput205, keyinput206, keyinput207;
  input keyinput208, keyinput209, keyinput210, keyinput211, keyinput212;
  input keyinput213, keyinput214, keyinput215, keyinput216, keyinput217;
  input keyinput218, keyinput219, keyinput220, keyinput221, keyinput222;
  input keyinput223, keyinput224, keyinput225, keyinput226, keyinput227;
  input keyinput228, keyinput229, keyinput230, keyinput231, keyinput232;
  input keyinput233, keyinput234, keyinput235, keyinput236, keyinput237;
  input keyinput238, keyinput239, keyinput240, keyinput241, keyinput242;
  input keyinput243, keyinput244, keyinput245, keyinput246, keyinput247;

  wire KeyWire_0_1 , KeyWire_0_2, keyinput_Wire_1;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31, keyinput32, keyinput33, keyinput34;
  input keyinput35, keyinput36, keyinput37, keyinput38, keyinput39;
  input keyinput40, keyinput41, keyinput42, keyinput43, keyinput44;
  input keyinput45, keyinput46, keyinput47, keyinput48, keyinput49;
  input keyinput50, keyinput51, keyinput52, keyinput53, keyinput54;
  input keyinput55, keyinput56, keyinput57, keyinput58, keyinput59;
  input keyinput60, keyinput61, keyinput62, keyinput63, keyinput64;
  input keyinput65, keyinput66, keyinput67, keyinput68, keyinput69;
  input keyinput70, keyinput71, keyinput72, keyinput73, keyinput74;
  input keyinput75, keyinput76, keyinput77, keyinput78, keyinput79;
  input keyinput80, keyinput81, keyinput82, keyinput83, keyinput84;
  input keyinput85, keyinput86, keyinput87, keyinput88, keyinput89;
  input keyinput90, keyinput91, keyinput92, keyinput93, keyinput94;
  input keyinput95, keyinput96, keyinput97, keyinput98, keyinput99;
  input keyinput100, keyinput101, keyinput102, keyinput103, keyinput104;
  input keyinput105, keyinput106, keyinput107, keyinput108, keyinput109;
  input keyinput110, keyinput111, keyinput112, keyinput113, keyinput114;
  input keyinput115, keyinput116, keyinput117, keyinput118, keyinput119;
  input keyinput120, keyinput121, keyinput122, keyinput123, keyinput124;
  input keyinput125, keyinput126, keyinput127;

  wire [0:127] keyinput_Wire_0;
  wire [0:65] KeyNOTWire_0;

input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;

output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;

wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877;

nand NAND4_1 (N269, N1, N8, N13, N17);
nand NAND4_2 (N270, N1, N26, N13, N17);
and AND3_3 (N273, N29, N36, N42);
and AND3_4 (N276, N1, N26, N51);
  nand NAND4_5 (keyinput_Wire_0[0], N1, N8, N51, N17);
  xnor keyGate_0_0(KeyNOTWire_0[0], keyinput0, keyinput_Wire_0[0]);
  not KeyNOTGate_0_0(N279, KeyNOTWire_0[0]);
nand NAND4_6 (N280, N1, N8, N13, N55);
nand NAND4_7 (N284, N59, N42, N68, N72);
nand NAND2_8 (N285, N29, N68);
nand NAND3_9 (N286, N59, N68, N74);
and AND3_10 (N287, N29, N75, N80);
  and AND3_11 (keyinput_Wire_0[1], N29, N75, N42);
  xor keyGate_0_1(N290, keyinput1, keyinput_Wire_0[1]);
and AND3_12 (N291, N29, N36, N80);
  and AND3_13 (keyinput_Wire_0[2], N29, N36, N42);
  xnor keyGate_0_2(KeyNOTWire_0[1], keyinput2, keyinput_Wire_0[2]);
  not KeyNOTGate_0_1(N292, KeyNOTWire_0[1]);
and AND3_14 (N293, N59, N75, N80);
and AND3_15 (N294, N59, N75, N42);
and AND3_16 (N295, N59, N36, N80);
and AND3_17 (N296, N59, N36, N42);
and AND2_18 (N297, N85, N86);
or OR2_19 (N298, N87, N88);
nand NAND2_20 (N301, N91, N96);
or OR2_21 (N302, N91, N96);
  nand NAND2_22 (keyinput_Wire_0[3], N101, N106);
  xor keyGate_0_3(N303, keyinput3, keyinput_Wire_0[3]);
  or OR2_23 (keyinput_Wire_0[4], N101, N106);
  xnor keyGate_0_4(KeyNOTWire_0[2], keyinput4, keyinput_Wire_0[4]);
  not KeyNOTGate_0_2(N304, KeyNOTWire_0[2]);
nand NAND2_24 (N305, N111, N116);
or OR2_25 (N306, N111, N116);
nand NAND2_26 (N307, N121, N126);
  or OR2_27 (keyinput_Wire_0[5], N121, N126);
  xor keyGate_0_5(KeyNOTWire_0[3], keyinput5, keyinput_Wire_0[5]);
  not KeyNOTGate_0_3(N308, KeyNOTWire_0[3]);
and AND2_28 (N309, N8, N138);
not NOT1_29 (N310, N268);
  and AND2_30 (keyinput_Wire_0[6], N51, N138);
  xor keyGate_0_6(N316, keyinput6, keyinput_Wire_0[6]);
and AND2_31 (N317, N17, N138);
  and AND2_32 (keyinput_Wire_0[7], N152, N138);
  xnor keyGate_0_7(KeyNOTWire_0[4], keyinput7, keyinput_Wire_0[7]);
  not KeyNOTGate_0_4(N318, KeyNOTWire_0[4]);
nand NAND2_33 (N319, N59, N156);
nor NOR2_34 (N322, N17, N42);
  and AND2_35 (keyinput_Wire_0[8], N17, N42);
  xor keyGate_0_8(KeyNOTWire_0[5], keyinput8, keyinput_Wire_0[8]);
  not KeyNOTGate_0_5(N323, KeyNOTWire_0[5]);
  nand NAND2_36 (keyinput_Wire_0[9], N159, N165);
  xnor keyGate_0_9(N324, keyinput9, keyinput_Wire_0[9]);
  or OR2_37 (keyinput_Wire_0[10], N159, N165);
  xor keyGate_0_10(KeyNOTWire_0[6], keyinput10, keyinput_Wire_0[10]);
  not KeyNOTGate_0_6(N325, KeyNOTWire_0[6]);
  nand NAND2_38 (keyinput_Wire_0[11], N171, N177);
  xnor keyGate_0_11(KeyNOTWire_0[7], keyinput11, keyinput_Wire_0[11]);
  not KeyNOTGate_0_7(N326, KeyNOTWire_0[7]);
  or OR2_39 (keyinput_Wire_0[12], N171, N177);
  xor keyGate_0_12(KeyNOTWire_0[8], keyinput12, keyinput_Wire_0[12]);
  not KeyNOTGate_0_8(N327, KeyNOTWire_0[8]);
nand NAND2_40 (N328, N183, N189);
  or OR2_41 (keyinput_Wire_0[13], N183, N189);
  xnor keyGate_0_13(N329, keyinput13, keyinput_Wire_0[13]);
nand NAND2_42 (N330, N195, N201);
  or OR2_43 (keyinput_Wire_0[14], N195, N201);
  xnor keyGate_0_14(N331, keyinput14, keyinput_Wire_0[14]);
  and AND2_44 (keyinput_Wire_0[15], N210, N91);
  xnor keyGate_0_15(KeyNOTWire_0[9], keyinput15, keyinput_Wire_0[15]);
  not KeyNOTGate_0_9(N332, KeyNOTWire_0[9]);
  and AND2_45 (keyinput_Wire_0[16], N210, N96);
  xor keyGate_0_16(KeyNOTWire_0[10], keyinput16, keyinput_Wire_0[16]);
  not KeyNOTGate_0_10(N333, KeyNOTWire_0[10]);
  and AND2_46 (keyinput_Wire_0[17], N210, N101);
  xor keyGate_0_17(KeyNOTWire_0[11], keyinput17, keyinput_Wire_0[17]);
  not KeyNOTGate_0_11(N334, KeyNOTWire_0[11]);
  and AND2_47 (keyinput_Wire_0[18], N210, N106);
  xnor keyGate_0_18(KeyNOTWire_0[12], keyinput18, keyinput_Wire_0[18]);
  not KeyNOTGate_0_12(N335, KeyNOTWire_0[12]);
and AND2_48 (N336, N210, N111);
and AND2_49 (N337, N255, N259);
and AND2_50 (N338, N210, N116);
and AND2_51 (N339, N255, N260);
  and AND2_52 (keyinput_Wire_0[19], N210, N121);
  xor keyGate_0_19(KeyNOTWire_0[13], keyinput19, keyinput_Wire_0[19]);
  not KeyNOTGate_0_13(N340, KeyNOTWire_0[13]);
  and AND2_53 (keyinput_Wire_0[20], N255, N267);
  xnor keyGate_0_20(N341, keyinput20, keyinput_Wire_0[20]);
not NOT1_54 (N342, N269);
not NOT1_55 (N343, N273);
or OR2_56 (N344, N270, N273);
  not NOT1_57 (keyinput_Wire_0[21], N276);
  xor keyGate_0_21(KeyNOTWire_0[14], keyinput21, keyinput_Wire_0[21]);
  not KeyNOTGate_0_14(N345, KeyNOTWire_0[14]);
  not NOT1_58 (keyinput_Wire_0[22], N276);
  xor keyGate_0_22(KeyNOTWire_0[15], keyinput22, keyinput_Wire_0[22]);
  not KeyNOTGate_0_15(N346, KeyNOTWire_0[15]);
not NOT1_59 (N347, N279);
nor NOR2_60 (N348, N280, N284);
or OR2_61 (N349, N280, N285);
or OR2_62 (N350, N280, N286);
not NOT1_63 (N351, N293);
not NOT1_64 (N352, N294);
not NOT1_65 (N353, N295);
not NOT1_66 (N354, N296);
nand NAND2_67 (N355, N89, N298);
and AND2_68 (N356, N90, N298);
nand NAND2_69 (N357, N301, N302);
  nand NAND2_70 (keyinput_Wire_0[23], N303, N304);
  xnor keyGate_0_23(KeyNOTWire_0[16], keyinput23, keyinput_Wire_0[23]);
  not KeyNOTGate_0_16(N360, KeyNOTWire_0[16]);
  nand NAND2_71 (keyinput_Wire_0[24], N305, N306);
  xnor keyGate_0_24(KeyNOTWire_0[17], keyinput24, keyinput_Wire_0[24]);
  not KeyNOTGate_0_17(N363, KeyNOTWire_0[17]);
nand NAND2_72 (N366, N307, N308);
not NOT1_73 (N369, N310);
nor NOR2_74 (N375, N322, N323);
  nand NAND2_75 (keyinput_Wire_0[25], N324, N325);
  xnor keyGate_0_25(N376, keyinput25, keyinput_Wire_0[25]);
  nand NAND2_76 (keyinput_Wire_0[26], N326, N327);
  xor keyGate_0_26(KeyNOTWire_0[18], keyinput26, keyinput_Wire_0[26]);
  not KeyNOTGate_0_18(N379, KeyNOTWire_0[18]);
  nand NAND2_77 (keyinput_Wire_0[27], N328, N329);
  xor keyGate_0_27(N382, keyinput27, keyinput_Wire_0[27]);
nand NAND2_78 (N385, N330, N331);
buf BUFF1_79 (N388, N290);
buf BUFF1_80 (N389, N291);
buf BUFF1_81 (N390, N292);
buf BUFF1_82 (N391, N297);
or OR2_83 (N392, N270, N343);
not NOT1_84 (N393, N345);
not NOT1_85 (N399, N346);
and AND2_86 (N400, N348, N73);
not NOT1_87 (N401, N349);
  not NOT1_88 (keyinput_Wire_0[28], N350);
  xnor keyGate_0_28(N402, keyinput28, keyinput_Wire_0[28]);
not NOT1_89 (N403, N355);
not NOT1_90 (N404, N357);
  not NOT1_91 (keyinput_Wire_0[29], N360);
  xor keyGate_0_29(KeyNOTWire_0[19], keyinput29, keyinput_Wire_0[29]);
  not KeyNOTGate_0_19(N405, KeyNOTWire_0[19]);
and AND2_92 (N406, N357, N360);
  not NOT1_93 (keyinput_Wire_0[30], N363);
  xnor keyGate_0_30(N407, keyinput30, keyinput_Wire_0[30]);
not NOT1_94 (N408, N366);
and AND2_95 (N409, N363, N366);
nand NAND2_96 (N410, N347, N352);
  not NOT1_97 (keyinput_Wire_0[31], N376);
  xnor keyGate_0_31(KeyNOTWire_0[20], keyinput31, keyinput_Wire_0[31]);
  not KeyNOTGate_0_20(N411, KeyNOTWire_0[20]);
  not NOT1_98 (keyinput_Wire_0[32], N379);
  xnor keyGate_0_32(N412, keyinput32, keyinput_Wire_0[32]);
and AND2_99 (N413, N376, N379);
not NOT1_100 (N414, N382);
  not NOT1_101 (keyinput_Wire_0[33], N385);
  xor keyGate_0_33(N415, keyinput33, keyinput_Wire_0[33]);
and AND2_102 (N416, N382, N385);
and AND2_103 (N417, N210, N369);
buf BUFF1_104 (N418, N342);
buf BUFF1_105 (N419, N344);
buf BUFF1_106 (N420, N351);
buf BUFF1_107 (N421, N353);
buf BUFF1_108 (N422, N354);
buf BUFF1_109 (N423, N356);
not NOT1_110 (N424, N400);
  and AND2_111 (keyinput_Wire_0[34], N404, N405);
  xnor keyGate_0_34(N425, keyinput34, keyinput_Wire_0[34]);
  and AND2_112 (keyinput_Wire_0[35], N407, N408);
  xnor keyGate_0_35(N426, keyinput35, keyinput_Wire_0[35]);
and AND3_113 (N427, N319, N393, N55);
and AND3_114 (N432, N393, N17, N287);
nand NAND3_115 (N437, N393, N287, N55);
  nand NAND4_116 (keyinput_Wire_0[36], N375, N59, N156, N393);
  xnor keyGate_0_36(KeyNOTWire_0[21], keyinput36, keyinput_Wire_0[36]);
  not KeyNOTGate_0_21(N442, KeyNOTWire_0[21]);
nand NAND3_117 (N443, N393, N319, N17);
  and AND2_118 (keyinput_Wire_0[37], N411, N412);
  xor keyGate_0_37(N444, keyinput37, keyinput_Wire_0[37]);
  and AND2_119 (keyinput_Wire_0[38], N414, N415);
  xnor keyGate_0_38(KeyNOTWire_0[22], keyinput38, keyinput_Wire_0[38]);
  not KeyNOTGate_0_22(N445, KeyNOTWire_0[22]);
buf BUFF1_120 (N446, N392);
buf BUFF1_121 (N447, N399);
buf BUFF1_122 (N448, N401);
buf BUFF1_123 (N449, N402);
buf BUFF1_124 (N450, N403);
  not NOT1_125 (keyinput_Wire_0[39], N424);
  xor keyGate_0_39(KeyNOTWire_0[23], keyinput39, keyinput_Wire_0[39]);
  not KeyNOTGate_0_23(N451, KeyNOTWire_0[23]);
nor NOR2_126 (N460, N406, N425);
  nor NOR2_127 (keyinput_Wire_0[40], N409, N426);
  xor keyGate_0_40(KeyNOTWire_0[24], keyinput40, keyinput_Wire_0[40]);
  not KeyNOTGate_0_24(N463, KeyNOTWire_0[24]);
  nand NAND2_128 (keyinput_Wire_0[41], N442, N410);
  xnor keyGate_0_41(N466, keyinput41, keyinput_Wire_0[41]);
  and AND2_129 (keyinput_Wire_0[42], N143, N427);
  xnor keyGate_0_42(N475, keyinput42, keyinput_Wire_0[42]);
  and AND2_130 (keyinput_Wire_0[43], N310, N432);
  xor keyGate_0_43(KeyNOTWire_0[25], keyinput43, keyinput_Wire_0[43]);
  not KeyNOTGate_0_25(N476, KeyNOTWire_0[25]);
and AND2_131 (N477, N146, N427);
and AND2_132 (N478, N310, N432);
  and AND2_133 (keyinput_Wire_0[44], N149, N427);
  xnor keyGate_0_44(KeyNOTWire_0[26], keyinput44, keyinput_Wire_0[44]);
  not KeyNOTGate_0_26(N479, KeyNOTWire_0[26]);
and AND2_134 (N480, N310, N432);
  and AND2_135 (keyinput_Wire_0[45], N153, N427);
  xnor keyGate_0_45(KeyNOTWire_0[27], keyinput45, keyinput_Wire_0[45]);
  not KeyNOTGate_0_27(N481, KeyNOTWire_0[27]);
  and AND2_136 (keyinput_Wire_0[46], N310, N432);
  xnor keyGate_0_46(KeyNOTWire_0[28], keyinput46, keyinput_Wire_0[46]);
  not KeyNOTGate_0_28(N482, KeyNOTWire_0[28]);
nand NAND2_137 (N483, N443, N1);
or OR2_138 (N488, N369, N437);
or OR2_139 (N489, N369, N437);
  or OR2_140 (keyinput_Wire_0[47], N369, N437);
  xor keyGate_0_47(N490, keyinput47, keyinput_Wire_0[47]);
  or OR2_141 (keyinput_Wire_0[48], N369, N437);
  xor keyGate_0_48(KeyNOTWire_0[29], keyinput48, keyinput_Wire_0[48]);
  not KeyNOTGate_0_29(N491, KeyNOTWire_0[29]);
nor NOR2_142 (N492, N413, N444);
  nor NOR2_143 (keyinput_Wire_0[49], N416, N445);
  xnor keyGate_0_49(KeyNOTWire_0[30], keyinput49, keyinput_Wire_0[49]);
  not KeyNOTGate_0_30(N495, KeyNOTWire_0[30]);
nand NAND2_144 (N498, N130, N460);
  or OR2_145 (keyinput_Wire_0[50], N130, N460);
  xnor keyGate_0_50(KeyNOTWire_0[31], keyinput50, keyinput_Wire_0[50]);
  not KeyNOTGate_0_31(N499, KeyNOTWire_0[31]);
  nand NAND2_146 (keyinput_Wire_0[51], N463, N135);
  xnor keyGate_0_51(KeyNOTWire_0[32], keyinput51, keyinput_Wire_0[51]);
  not KeyNOTGate_0_32(N500, KeyNOTWire_0[32]);
or OR2_147 (N501, N463, N135);
and AND2_148 (N502, N91, N466);
nor NOR2_149 (N503, N475, N476);
and AND2_150 (N504, N96, N466);
nor NOR2_151 (N505, N477, N478);
and AND2_152 (N506, N101, N466);
  nor NOR2_153 (keyinput_Wire_0[52], N479, N480);
  xor keyGate_0_52(KeyNOTWire_0[33], keyinput52, keyinput_Wire_0[52]);
  not KeyNOTGate_0_33(N507, KeyNOTWire_0[33]);
and AND2_154 (N508, N106, N466);
nor NOR2_155 (N509, N481, N482);
and AND2_156 (N510, N143, N483);
  and AND2_157 (keyinput_Wire_0[53], N111, N466);
  xor keyGate_0_53(N511, keyinput53, keyinput_Wire_0[53]);
and AND2_158 (N512, N146, N483);
and AND2_159 (N513, N116, N466);
and AND2_160 (N514, N149, N483);
  and AND2_161 (keyinput_Wire_0[54], N121, N466);
  xor keyGate_0_54(KeyNOTWire_0[34], keyinput54, keyinput_Wire_0[54]);
  not KeyNOTGate_0_34(N515, KeyNOTWire_0[34]);
and AND2_162 (N516, N153, N483);
and AND2_163 (N517, N126, N466);
  nand NAND2_164 (keyinput_Wire_0[55], N130, N492);
  xnor keyGate_0_55(KeyNOTWire_0[35], keyinput55, keyinput_Wire_0[55]);
  not KeyNOTGate_0_35(N518, KeyNOTWire_0[35]);
  or OR2_165 (keyinput_Wire_0[56], N130, N492);
  xnor keyGate_0_56(KeyNOTWire_0[36], keyinput56, keyinput_Wire_0[56]);
  not KeyNOTGate_0_36(N519, KeyNOTWire_0[36]);
nand NAND2_166 (N520, N495, N207);
or OR2_167 (N521, N495, N207);
  and AND2_168 (keyinput_Wire_0[57], N451, N159);
  xnor keyGate_0_57(KeyNOTWire_0[37], keyinput57, keyinput_Wire_0[57]);
  not KeyNOTGate_0_37(N522, KeyNOTWire_0[37]);
and AND2_169 (N523, N451, N165);
and AND2_170 (N524, N451, N171);
and AND2_171 (N525, N451, N177);
and AND2_172 (N526, N451, N183);
nand NAND2_173 (N527, N451, N189);
nand NAND2_174 (N528, N451, N195);
nand NAND2_175 (N529, N451, N201);
nand NAND2_176 (N530, N498, N499);
nand NAND2_177 (N533, N500, N501);
  nor NOR2_178 (keyinput_Wire_0[58], N309, N502);
  xnor keyGate_0_58(N536, keyinput58, keyinput_Wire_0[58]);
nor NOR2_179 (N537, N316, N504);
nor NOR2_180 (N538, N317, N506);
nor NOR2_181 (N539, N318, N508);
nor NOR2_182 (N540, N510, N511);
  nor NOR2_183 (keyinput_Wire_0[59], N512, N513);
  xor keyGate_0_59(KeyNOTWire_0[38], keyinput59, keyinput_Wire_0[59]);
  not KeyNOTGate_0_38(N541, KeyNOTWire_0[38]);
  nor NOR2_184 (keyinput_Wire_0[60], N514, N515);
  xnor keyGate_0_60(N542, keyinput60, keyinput_Wire_0[60]);
nor NOR2_185 (N543, N516, N517);
nand NAND2_186 (N544, N518, N519);
nand NAND2_187 (N547, N520, N521);
not NOT1_188 (N550, N530);
not NOT1_189 (N551, N533);
and AND2_190 (N552, N530, N533);
nand NAND2_191 (N553, N536, N503);
nand NAND2_192 (N557, N537, N505);
  nand NAND2_193 (keyinput_Wire_0[61], N538, N507);
  xnor keyGate_0_61(KeyNOTWire_0[39], keyinput61, keyinput_Wire_0[61]);
  not KeyNOTGate_0_39(N561, KeyNOTWire_0[39]);
nand NAND2_194 (N565, N539, N509);
nand NAND2_195 (N569, N488, N540);
  nand NAND2_196 (keyinput_Wire_0[62], N489, N541);
  xor keyGate_0_62(KeyNOTWire_0[40], keyinput62, keyinput_Wire_0[62]);
  not KeyNOTGate_0_40(N573, KeyNOTWire_0[40]);
nand NAND2_197 (N577, N490, N542);
nand NAND2_198 (N581, N491, N543);
not NOT1_199 (N585, N544);
not NOT1_200 (N586, N547);
  and AND2_201 (keyinput_Wire_0[63], N544, N547);
  xor keyGate_0_63(N587, keyinput63, keyinput_Wire_0[63]);
and AND2_202 (N588, N550, N551);
  and AND2_203 (keyinput_Wire_0[64], N585, N586);
  xnor keyGate_0_64(N589, keyinput64, keyinput_Wire_0[64]);
nand NAND2_204 (N590, N553, N159);
or OR2_205 (N593, N553, N159);
and AND2_206 (N596, N246, N553);
nand NAND2_207 (N597, N557, N165);
  or OR2_208 (keyinput_Wire_0[65], N557, N165);
  xnor keyGate_0_65(KeyNOTWire_0[41], keyinput65, keyinput_Wire_0[65]);
  not KeyNOTGate_0_41(N600, KeyNOTWire_0[41]);
  and AND2_209 (keyinput_Wire_0[66], N246, N557);
  xor keyGate_0_66(N605, keyinput66, keyinput_Wire_0[66]);
nand NAND2_210 (N606, N561, N171);
  or OR2_211 (keyinput_Wire_0[67], N561, N171);
  xor keyGate_0_67(N609, keyinput67, keyinput_Wire_0[67]);
and AND2_212 (N615, N246, N561);
nand NAND2_213 (N616, N565, N177);
or OR2_214 (N619, N565, N177);
and AND2_215 (N624, N246, N565);
nand NAND2_216 (N625, N569, N183);
or OR2_217 (N628, N569, N183);
  and AND2_218 (keyinput_Wire_0[68], N246, N569);
  xor keyGate_0_68(KeyNOTWire_0[42], keyinput68, keyinput_Wire_0[68]);
  not KeyNOTGate_0_42(N631, KeyNOTWire_0[42]);
nand NAND2_219 (N632, N573, N189);
  or OR2_220 (keyinput_Wire_0[69], N573, N189);
  xor keyGate_0_69(N635, keyinput69, keyinput_Wire_0[69]);
and AND2_221 (N640, N246, N573);
nand NAND2_222 (N641, N577, N195);
or OR2_223 (N644, N577, N195);
and AND2_224 (N650, N246, N577);
nand NAND2_225 (N651, N581, N201);
  or OR2_226 (keyinput_Wire_0[70], N581, N201);
  xor keyGate_0_70(KeyNOTWire_0[43], keyinput70, keyinput_Wire_0[70]);
  not KeyNOTGate_0_43(N654, KeyNOTWire_0[43]);
and AND2_227 (N659, N246, N581);
  nor NOR2_228 (keyinput_Wire_0[71], N552, N588);
  xnor keyGate_0_71(N660, keyinput71, keyinput_Wire_0[71]);
nor NOR2_229 (N661, N587, N589);
  not NOT1_230 (keyinput_Wire_0[72], N590);
  xor keyGate_0_72(N662, keyinput72, keyinput_Wire_0[72]);
and AND2_231 (N665, N593, N590);
  nor NOR2_232 (keyinput_Wire_0[73], N596, N522);
  xnor keyGate_0_73(KeyNOTWire_0[44], keyinput73, keyinput_Wire_0[73]);
  not KeyNOTGate_0_44(N669, KeyNOTWire_0[44]);
not NOT1_233 (N670, N597);
and AND2_234 (N673, N600, N597);
nor NOR2_235 (N677, N605, N523);
  not NOT1_236 (keyinput_Wire_0[74], N606);
  xnor keyGate_0_74(KeyNOTWire_0[45], keyinput74, keyinput_Wire_0[74]);
  not KeyNOTGate_0_45(N678, KeyNOTWire_0[45]);
  and AND2_237 (keyinput_Wire_0[75], N609, N606);
  xnor keyGate_0_75(N682, keyinput75, keyinput_Wire_0[75]);
  nor NOR2_238 (keyinput_Wire_0[76], N615, N524);
  xor keyGate_0_76(N686, keyinput76, keyinput_Wire_0[76]);
  not NOT1_239 (keyinput_Wire_0[77], N616);
  xnor keyGate_0_77(KeyNOTWire_0[46], keyinput77, keyinput_Wire_0[77]);
  not KeyNOTGate_0_46(N687, KeyNOTWire_0[46]);
  and AND2_240 (keyinput_Wire_0[78], N619, N616);
  xnor keyGate_0_78(KeyNOTWire_0[47], keyinput78, keyinput_Wire_0[78]);
  not KeyNOTGate_0_47(N692, KeyNOTWire_0[47]);
  nor NOR2_241 (keyinput_Wire_0[79], N624, N525);
  xnor keyGate_0_79(N696, keyinput79, keyinput_Wire_0[79]);
not NOT1_242 (N697, N625);
  and AND2_243 (keyinput_Wire_0[80], N628, N625);
  xor keyGate_0_80(N700, keyinput80, keyinput_Wire_0[80]);
nor NOR2_244 (N704, N631, N526);
not NOT1_245 (N705, N632);
  and AND2_246 (keyinput_Wire_0[81], N635, N632);
  xnor keyGate_0_81(N708, keyinput81, keyinput_Wire_0[81]);
nor NOR2_247 (N712, N337, N640);
not NOT1_248 (N713, N641);
and AND2_249 (N717, N644, N641);
nor NOR2_250 (N721, N339, N650);
not NOT1_251 (N722, N651);
  and AND2_252 (keyinput_Wire_0[82], N654, N651);
  xnor keyGate_0_82(N727, keyinput82, keyinput_Wire_0[82]);
nor NOR2_253 (N731, N341, N659);
nand NAND2_254 (N732, N654, N261);
nand NAND3_255 (N733, N644, N654, N261);
  nand NAND4_256 (keyinput_Wire_0[83], N635, N644, N654, N261);
  xnor keyGate_0_83(N734, keyinput83, keyinput_Wire_0[83]);
  not NOT1_257 (keyinput_Wire_0[84], N662);
  xor keyGate_0_84(N735, keyinput84, keyinput_Wire_0[84]);
  and AND2_258 (keyinput_Wire_0[85], N228, N665);
  xnor keyGate_0_85(N736, keyinput85, keyinput_Wire_0[85]);
  and AND2_259 (keyinput_Wire_0[86], N237, N662);
  xnor keyGate_0_86(KeyNOTWire_0[48], keyinput86, keyinput_Wire_0[86]);
  not KeyNOTGate_0_48(N737, KeyNOTWire_0[48]);
not NOT1_260 (N738, N670);
and AND2_261 (N739, N228, N673);
  and AND2_262 (keyinput_Wire_0[87], N237, N670);
  xnor keyGate_0_87(KeyNOTWire_0[49], keyinput87, keyinput_Wire_0[87]);
  not KeyNOTGate_0_49(N740, KeyNOTWire_0[49]);
not NOT1_263 (N741, N678);
  and AND2_264 (keyinput_Wire_0[88], N228, N682);
  xnor keyGate_0_88(N742, keyinput88, keyinput_Wire_0[88]);
  and AND2_265 (keyinput_Wire_0[89], N237, N678);
  xnor keyGate_0_89(N743, keyinput89, keyinput_Wire_0[89]);
not NOT1_266 (N744, N687);
and AND2_267 (N745, N228, N692);
and AND2_268 (N746, N237, N687);
not NOT1_269 (N747, N697);
and AND2_270 (N748, N228, N700);
and AND2_271 (N749, N237, N697);
not NOT1_272 (N750, N705);
and AND2_273 (N751, N228, N708);
and AND2_274 (N752, N237, N705);
  not NOT1_275 (keyinput_Wire_0[90], N713);
  xnor keyGate_0_90(N753, keyinput90, keyinput_Wire_0[90]);
and AND2_276 (N754, N228, N717);
  and AND2_277 (keyinput_Wire_0[91], N237, N713);
  xnor keyGate_0_91(N755, keyinput91, keyinput_Wire_0[91]);
not NOT1_278 (N756, N722);
nor NOR2_279 (N757, N727, N261);
and AND2_280 (N758, N727, N261);
and AND2_281 (N759, N228, N727);
and AND2_282 (N760, N237, N722);
  nand NAND2_283 (keyinput_Wire_0[92], N644, N722);
  xor keyGate_0_92(N761, keyinput92, keyinput_Wire_0[92]);
nand NAND2_284 (N762, N635, N713);
  nand NAND3_285 (keyinput_Wire_0[93], N635, N644, N722);
  xor keyGate_0_93(N763, keyinput93, keyinput_Wire_0[93]);
nand NAND2_286 (N764, N609, N687);
  nand NAND2_287 (keyinput_Wire_0[94], N600, N678);
  xnor keyGate_0_94(KeyNOTWire_0[50], keyinput94, keyinput_Wire_0[94]);
  not KeyNOTGate_0_50(N765, KeyNOTWire_0[50]);
  nand NAND3_288 (keyinput_Wire_0[95], N600, N609, N687);
  xor keyGate_0_95(N766, keyinput95, keyinput_Wire_0[95]);
buf BUFF1_289 (N767, N660);
  buf BUFF1_290 (keyinput_Wire_1, N661);
  xor keyGate_1_5(N768, KeyWire_0_2, keyinput_Wire_1);
nor NOR2_291 (N769, N736, N737);
  nor NOR2_292 (keyinput_Wire_0[96], N739, N740);
  xnor keyGate_0_96(N770, keyinput96, keyinput_Wire_0[96]);
nor NOR2_293 (N771, N742, N743);
  nor NOR2_294 (keyinput_Wire_0[97], N745, N746);
  xnor keyGate_0_97(KeyNOTWire_0[51], keyinput97, keyinput_Wire_0[97]);
  not KeyNOTGate_0_51(N772, KeyNOTWire_0[51]);
  nand NAND4_295 (keyinput_Wire_0[98], N750, N762, N763, N734);
  xor keyGate_0_98(N773, keyinput98, keyinput_Wire_0[98]);
nor NOR2_296 (N777, N748, N749);
nand NAND3_297 (N778, N753, N761, N733);
  nor NOR2_298 (keyinput_Wire_0[99], N751, N752);
  xor keyGate_0_99(KeyNOTWire_0[52], keyinput99, keyinput_Wire_0[99]);
  not KeyNOTGate_0_52(N781, KeyNOTWire_0[52]);
nand NAND2_299 (N782, N756, N732);
nor NOR2_300 (N785, N754, N755);
nor NOR2_301 (N786, N757, N758);
nor NOR2_302 (N787, N759, N760);
  nor NOR2_303 (keyinput_Wire_0[100], N700, N773);
  xnor keyGate_0_100(KeyNOTWire_0[53], keyinput100, keyinput_Wire_0[100]);
  not KeyNOTGate_0_53(N788, KeyNOTWire_0[53]);
and AND2_304 (N789, N700, N773);
nor NOR2_305 (N790, N708, N778);
  and AND2_306 (keyinput_Wire_0[101], N708, N778);
  xnor keyGate_0_101(N791, keyinput101, keyinput_Wire_0[101]);
  nor NOR2_307 (keyinput_Wire_0[102], N717, N782);
  xnor keyGate_0_102(N792, keyinput102, keyinput_Wire_0[102]);
  and AND2_308 (keyinput_Wire_0[103], N717, N782);
  xor keyGate_0_103(KeyNOTWire_0[54], keyinput103, keyinput_Wire_0[103]);
  not KeyNOTGate_0_54(N793, KeyNOTWire_0[54]);
and AND2_309 (N794, N219, N786);
  nand NAND2_310 (keyinput_Wire_0[104], N628, N773);
  xor keyGate_0_104(N795, keyinput104, keyinput_Wire_0[104]);
nand NAND2_311 (N796, N795, N747);
nor NOR2_312 (N802, N788, N789);
nor NOR2_313 (N803, N790, N791);
nor NOR2_314 (N804, N792, N793);
nor NOR2_315 (N805, N340, N794);
nor NOR2_316 (N806, N692, N796);
and AND2_317 (N807, N692, N796);
  and AND2_318 (keyinput_Wire_0[105], N219, N802);
  xnor keyGate_0_105(N808, keyinput105, keyinput_Wire_0[105]);
and AND2_319 (N809, N219, N803);
  and AND2_320 (keyinput_Wire_0[106], N219, N804);
  xor keyGate_0_106(KeyNOTWire_0[55], keyinput106, keyinput_Wire_0[106]);
  not KeyNOTGate_0_55(N810, KeyNOTWire_0[55]);
  nand NAND4_321 (keyinput_Wire_0[107], N805, N787, N731, N529);
  xor keyGate_0_107(N811, keyinput107, keyinput_Wire_0[107]);
  nand NAND2_322 (keyinput_Wire_0[108], N619, N796);
  xnor keyGate_0_108(KeyNOTWire_0[56], keyinput108, keyinput_Wire_0[108]);
  not KeyNOTGate_0_56(N812, KeyNOTWire_0[56]);
nand NAND3_323 (N813, N609, N619, N796);
nand NAND4_324 (N814, N600, N609, N619, N796);
nand NAND4_325 (N815, N738, N765, N766, N814);
nand NAND3_326 (N819, N741, N764, N813);
nand NAND2_327 (N822, N744, N812);
  nor NOR2_328 (keyinput_Wire_0[109], N806, N807);
  xor keyGate_0_109(N825, keyinput109, keyinput_Wire_0[109]);
nor NOR2_329 (N826, N335, N808);
nor NOR2_330 (N827, N336, N809);
nor NOR2_331 (N828, N338, N810);
  not NOT1_332 (keyinput_Wire_0[110], N811);
  xor keyGate_0_110(N829, keyinput110, keyinput_Wire_0[110]);
  nor NOR2_333 (keyinput_Wire_0[111], N665, N815);
  xor keyGate_0_111(KeyNOTWire_0[57], keyinput111, keyinput_Wire_0[111]);
  not KeyNOTGate_0_57(N830, KeyNOTWire_0[57]);
and AND2_334 (N831, N665, N815);
nor NOR2_335 (N832, N673, N819);
and AND2_336 (N833, N673, N819);
  nor NOR2_337 (keyinput_Wire_0[112], N682, N822);
  xor keyGate_0_112(KeyNOTWire_0[58], keyinput112, keyinput_Wire_0[112]);
  not KeyNOTGate_0_58(N834, KeyNOTWire_0[58]);
  and AND2_338 (keyinput_Wire_0[113], N682, N822);
  xnor keyGate_0_113(N835, keyinput113, keyinput_Wire_0[113]);
and AND2_339 (N836, N219, N825);
  nand NAND3_340 (keyinput_Wire_0[114], N826, N777, N704);
  xnor keyGate_0_114(KeyNOTWire_0[59], keyinput114, keyinput_Wire_0[114]);
  not KeyNOTGate_0_59(N837, KeyNOTWire_0[59]);
  nand NAND4_341 (keyinput_Wire_0[115], N827, N781, N712, N527);
  xnor keyGate_0_115(KeyNOTWire_0[60], keyinput115, keyinput_Wire_0[115]);
  not KeyNOTGate_0_60(N838, KeyNOTWire_0[60]);
nand NAND4_342 (N839, N828, N785, N721, N528);
not NOT1_343 (N840, N829);
nand NAND2_344 (N841, N815, N593);
  nor NOR2_345 (keyinput_Wire_0[116], N830, N831);
  xor keyGate_0_116(N842, keyinput116, keyinput_Wire_0[116]);
nor NOR2_346 (N843, N832, N833);
nor NOR2_347 (N844, N834, N835);
nor NOR2_348 (N845, N334, N836);
not NOT1_349 (N846, N837);
not NOT1_350 (N847, N838);
not NOT1_351 (N848, N839);
  and AND2_352 (keyinput_Wire_0[117], N735, N841);
  xnor keyGate_0_117(N849, keyinput117, keyinput_Wire_0[117]);
buf BUFF1_353 (N850, N840);
  and AND2_354 (keyinput_Wire_0[118], N219, N842);
  xnor keyGate_0_118(N851, keyinput118, keyinput_Wire_0[118]);
and AND2_355 (N852, N219, N843);
  and AND2_356 (keyinput_Wire_0[119], N219, N844);
  xnor keyGate_0_119(KeyNOTWire_0[61], keyinput119, keyinput_Wire_0[119]);
  not KeyNOTGate_0_61(N853, KeyNOTWire_0[61]);
nand NAND3_357 (N854, N845, N772, N696);
  not NOT1_358 (keyinput_Wire_0[120], N846);
  xnor keyGate_0_120(N855, keyinput120, keyinput_Wire_0[120]);
  not NOT1_359 (keyinput_Wire_0[121], N847);
  xor keyGate_0_121(KeyNOTWire_0[62], keyinput121, keyinput_Wire_0[121]);
  not KeyNOTGate_0_62(N856, KeyNOTWire_0[62]);
  not NOT1_360 (keyinput_Wire_0[122], N848);
  xnor keyGate_0_122(N857, keyinput122, keyinput_Wire_0[122]);
not NOT1_361 (N858, N849);
nor NOR2_362 (N859, N417, N851);
nor NOR2_363 (N860, N332, N852);
nor NOR2_364 (N861, N333, N853);
  not NOT1_365 (keyinput_Wire_0[123], N854);
  xnor keyGate_0_123(KeyNOTWire_0[63], keyinput123, keyinput_Wire_0[123]);
  not KeyNOTGate_0_63(N862, KeyNOTWire_0[63]);
buf BUFF1_366 (KeyWire_0_1, N855);
  xor flip_it (N863, KeyWire_0_1, KeyWire_0_2 );
buf BUFF1_367 (N864, N856);
buf BUFF1_368 (N865, N857);
buf BUFF1_369 (N866, N858);
nand NAND3_370 (N867, N859, N769, N669);
nand NAND3_371 (N868, N860, N770, N677);
nand NAND3_372 (N869, N861, N771, N686);
  not NOT1_373 (keyinput_Wire_0[124], N862);
  xnor keyGate_0_124(KeyNOTWire_0[64], keyinput124, keyinput_Wire_0[124]);
  not KeyNOTGate_0_64(N870, KeyNOTWire_0[64]);
not NOT1_374 (N871, N867);
not NOT1_375 (N872, N868);
  not NOT1_376 (keyinput_Wire_0[125], N869);
  xor keyGate_0_125(N873, keyinput125, keyinput_Wire_0[125]);
buf BUFF1_377 (N874, N870);
  not NOT1_378 (keyinput_Wire_0[126], N871);
  xnor keyGate_0_126(N875, keyinput126, keyinput_Wire_0[126]);
not NOT1_379 (N876, N872);
  not NOT1_380 (keyinput_Wire_0[127], N873);
  xor keyGate_0_127(KeyNOTWire_0[65], keyinput127, keyinput_Wire_0[127]);
  not KeyNOTGate_0_65(N877, KeyNOTWire_0[65]);
buf BUFF1_381 (N878, N875);
buf BUFF1_382 (N879, N876);
buf BUFF1_383 (N880, N877);

AntiSAT some_name( KeyWire_0_2, N59, N126, N183, N165, N156, N237, N8, N138, N207, N1, N91, N246, N68, N26, N135, N90, N261, N121, N177, N268, N130, N85, N195, N36, N74, N96, N159, N111, N267, N219, N13, N73, N116, N143, N260, N72, N75, N152, N86, N201, N89, N149, N228, N80, N55, N259, N101, N189, N42, N106, N88, N153, N17, N146, N87, N51, N29, N255, N210, N171, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, keyinput245, keyinput246, keyinput247,
       keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
       keyinput253, keyinput254, keyinput255, keyinput256, keyinput257,
       keyinput258, keyinput259, keyinput260, keyinput261, keyinput262,
       keyinput263, keyinput264, keyinput265, keyinput266, keyinput267,
       keyinput268, keyinput269, keyinput270, keyinput271, keyinput272,
       keyinput273, keyinput274, keyinput275, keyinput276, keyinput277,
       keyinput278, keyinput279, keyinput280, keyinput281, keyinput282,
       keyinput283, keyinput284, keyinput285, keyinput286, keyinput287,
       keyinput288, keyinput289, keyinput290, keyinput291, keyinput292,
       keyinput293, keyinput294, keyinput295, keyinput296, keyinput297,
       keyinput298, keyinput299, keyinput300, keyinput301, keyinput302,
       keyinput303, keyinput304, keyinput305, keyinput306, keyinput307);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N59, N126, N183, N165, N156, N237, N8, N138, N207, N1, N91, N246, N68, N26, N135, N90, N261, N121, N177, N268, N130, N85, N195, N36, N74, N96, N159, N111, N267, N219, N13, N73, N116, N143, N260, N72, N75, N152, N86, N201, N89, N149, N228, N80, N55, N259, N101, N189, N42, N106, N88, N153, N17, N146, N87, N51, N29, N255, N210, N171, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, keyinput245, keyinput246, keyinput247 ,
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
        keyinput253, keyinput254, keyinput255, keyinput256, keyinput257,
        keyinput258, keyinput259, keyinput260, keyinput261, keyinput262,
        keyinput263, keyinput264, keyinput265, keyinput266, keyinput267,
        keyinput268, keyinput269, keyinput270, keyinput271, keyinput272,
        keyinput273, keyinput274, keyinput275, keyinput276, keyinput277,
        keyinput278, keyinput279, keyinput280, keyinput281, keyinput282,
        keyinput283, keyinput284, keyinput285, keyinput286, keyinput287,
        keyinput288, keyinput289, keyinput290, keyinput291, keyinput292,
        keyinput293, keyinput294, keyinput295, keyinput296, keyinput297,
        keyinput298, keyinput299, keyinput300, keyinput301, keyinput302,
        keyinput303, keyinput304, keyinput305, keyinput306, keyinput307);

  input keyinput248, keyinput249, keyinput250, keyinput251, keyinput252;
  input keyinput253, keyinput254, keyinput255, keyinput256, keyinput257;
  input keyinput258, keyinput259, keyinput260, keyinput261, keyinput262;
  input keyinput263, keyinput264, keyinput265, keyinput266, keyinput267;
  input keyinput268, keyinput269, keyinput270, keyinput271, keyinput272;
  input keyinput273, keyinput274, keyinput275, keyinput276, keyinput277;
  input keyinput278, keyinput279, keyinput280, keyinput281, keyinput282;
  input keyinput283, keyinput284, keyinput285, keyinput286, keyinput287;
  input keyinput288, keyinput289, keyinput290, keyinput291, keyinput292;
  input keyinput293, keyinput294, keyinput295, keyinput296, keyinput297;
  input keyinput298, keyinput299, keyinput300, keyinput301, keyinput302;
  input keyinput303, keyinput304, keyinput305, keyinput306, keyinput307;

  wire [0:59] keyNTin_Wire_1;
  wire [0:26] KeyNOTWire_1;

  input N59, N126, N183, N165, N156, N237, N8, N138, N207, N1, N91, N246, N68, N26, N135, N90, N261, N121, N177, N268, N130, N85, N195, N36, N74, N96, N159, N111, N267, N219, N13, N73, N116, N143, N260, N72, N75, N152, N86, N201, N89, N149, N228, N80, N55, N259, N101, N189, N42, N106, N88, N153, N17, N146, N87, N51, N29, N255, N210, N171;
  input keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, keyinput245, keyinput246, keyinput247;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83, newWire_84, newWire_85, newWire_86, newWire_87, newWire_88, newWire_89, newWire_90, newWire_91, newWire_92, newWire_93, newWire_94, newWire_95, newWire_96, newWire_97, newWire_98, newWire_99, newWire_100, newWire_101, newWire_102, newWire_103, newWire_104, newWire_105, newWire_106, newWire_107, newWire_108, newWire_109, newWire_110, newWire_111, newWire_112, newWire_113, newWire_114, newWire_115, newWire_116, newWire_117, newWire_118, newWire_119, newWire_120, newWire_121 ;

  xnor KeyGate0 (keyNTin_Wire_1[0], N59, keyinput128);
  xor keyNTinGate_1_0(KeyNOTWire_1[0], keyinput248, keyNTin_Wire_1[0]);
  not KeyNOTGate_1_0(newWire_0, KeyNOTWire_1[0]);
  xnor KeyGate1 (newWire_1, N126, keyinput129);
  xor  KeyGate2 (keyNTin_Wire_1[1], N183, keyinput130);
  xnor keyNTinGate_1_1(newWire_2, keyinput249, keyNTin_Wire_1[1]);
  xor  KeyGate3 (newWire_3, N165, keyinput131);
  xnor KeyGate4 (keyNTin_Wire_1[2], N156, keyinput132);
  xnor keyNTinGate_1_2(newWire_4, keyinput250, keyNTin_Wire_1[2]);
  xor  KeyGate5 (newWire_5, N237, keyinput133);
  xor  KeyGate6 (keyNTin_Wire_1[3], N8, keyinput134);
  xnor keyNTinGate_1_3(newWire_6, keyinput251, keyNTin_Wire_1[3]);
  xor  KeyGate7 (keyNTin_Wire_1[4], N138, keyinput135);
  xor keyNTinGate_1_4(KeyNOTWire_1[1], keyinput252, keyNTin_Wire_1[4]);
  not KeyNOTGate_1_1(newWire_7, KeyNOTWire_1[1]);
  xnor KeyGate8 (newWire_8, N207, keyinput136);
  xnor KeyGate9 (newWire_9, N1, keyinput137);
  xnor KeyGate10 (newWire_10, N91, keyinput138);
  xnor KeyGate11 (keyNTin_Wire_1[5], N246, keyinput139);
  xnor keyNTinGate_1_5(newWire_11, keyinput253, keyNTin_Wire_1[5]);
  xnor KeyGate12 (keyNTin_Wire_1[6], N68, keyinput140);
  xnor keyNTinGate_1_6(newWire_12, keyinput254, keyNTin_Wire_1[6]);
  xor  KeyGate13 (keyNTin_Wire_1[7], N26, keyinput141);
  xor keyNTinGate_1_7(KeyNOTWire_1[2], keyinput255, keyNTin_Wire_1[7]);
  not KeyNOTGate_1_2(newWire_13, KeyNOTWire_1[2]);
  xnor KeyGate14 (newWire_14, N135, keyinput142);
  xnor KeyGate15 (newWire_15, N90, keyinput143);
  xor  KeyGate16 (keyNTin_Wire_1[8], N261, keyinput144);
  xor keyNTinGate_1_8(KeyNOTWire_1[3], keyinput256, keyNTin_Wire_1[8]);
  not KeyNOTGate_1_3(newWire_16, KeyNOTWire_1[3]);
  xor  KeyGate17 (newWire_17, N121, keyinput145);
  xnor KeyGate18 (keyNTin_Wire_1[9], N177, keyinput146);
  xnor keyNTinGate_1_9(newWire_18, keyinput257, keyNTin_Wire_1[9]);
  xnor KeyGate19 (keyNTin_Wire_1[10], N268, keyinput147);
  xnor keyNTinGate_1_10(newWire_19, keyinput258, keyNTin_Wire_1[10]);
  xnor KeyGate20 (keyNTin_Wire_1[11], N130, keyinput148);
  xnor keyNTinGate_1_11(KeyNOTWire_1[4], keyinput259, keyNTin_Wire_1[11]);
  not KeyNOTGate_1_4(newWire_20, KeyNOTWire_1[4]);
  xnor KeyGate21 (newWire_21, N85, keyinput149);
  xor  KeyGate22 (newWire_22, N195, keyinput150);
  xnor KeyGate23 (newWire_23, N36, keyinput151);
  xnor KeyGate24 (keyNTin_Wire_1[12], N74, keyinput152);
  xnor keyNTinGate_1_12(newWire_24, keyinput260, keyNTin_Wire_1[12]);
  xor  KeyGate25 (keyNTin_Wire_1[13], N96, keyinput153);
  xnor keyNTinGate_1_13(KeyNOTWire_1[5], keyinput261, keyNTin_Wire_1[13]);
  not KeyNOTGate_1_5(newWire_25, KeyNOTWire_1[5]);
  xnor KeyGate26 (keyNTin_Wire_1[14], N159, keyinput154);
  xor keyNTinGate_1_14(newWire_26, keyinput262, keyNTin_Wire_1[14]);
  xnor KeyGate27 (newWire_27, N111, keyinput155);
  xor  KeyGate28 (newWire_28, N267, keyinput156);
  xnor KeyGate29 (newWire_29, N219, keyinput157);
  xnor KeyGate30 (keyNTin_Wire_1[15], N13, keyinput158);
  xnor keyNTinGate_1_15(newWire_30, keyinput263, keyNTin_Wire_1[15]);
  xnor KeyGate31 (keyNTin_Wire_1[16], N73, keyinput159);
  xnor keyNTinGate_1_16(KeyNOTWire_1[6], keyinput264, keyNTin_Wire_1[16]);
  not KeyNOTGate_1_6(newWire_31, KeyNOTWire_1[6]);
  xor  KeyGate32 (newWire_32, N116, keyinput160);
  xor  KeyGate33 (newWire_33, N143, keyinput161);
  xnor KeyGate34 (newWire_34, N260, keyinput162);
  xor  KeyGate35 (keyNTin_Wire_1[17], N72, keyinput163);
  xnor keyNTinGate_1_17(KeyNOTWire_1[7], keyinput265, keyNTin_Wire_1[17]);
  not KeyNOTGate_1_7(newWire_35, KeyNOTWire_1[7]);
  xnor KeyGate36 (keyNTin_Wire_1[18], N75, keyinput164);
  xor keyNTinGate_1_18(newWire_36, keyinput266, keyNTin_Wire_1[18]);
  xor  KeyGate37 (keyNTin_Wire_1[19], N152, keyinput165);
  xnor keyNTinGate_1_19(KeyNOTWire_1[8], keyinput267, keyNTin_Wire_1[19]);
  not KeyNOTGate_1_8(newWire_37, KeyNOTWire_1[8]);
  xor  KeyGate38 (newWire_38, N86, keyinput166);
  xor  KeyGate39 (keyNTin_Wire_1[20], N201, keyinput167);
  xnor keyNTinGate_1_20(newWire_39, keyinput268, keyNTin_Wire_1[20]);
  xnor KeyGate40 (keyNTin_Wire_1[21], N89, keyinput168);
  xnor keyNTinGate_1_21(KeyNOTWire_1[9], keyinput269, keyNTin_Wire_1[21]);
  not KeyNOTGate_1_9(newWire_40, KeyNOTWire_1[9]);
  xnor KeyGate41 (keyNTin_Wire_1[22], N149, keyinput169);
  xor keyNTinGate_1_22(newWire_41, keyinput270, keyNTin_Wire_1[22]);
  xnor KeyGate42 (newWire_42, N228, keyinput170);
  xnor KeyGate43 (newWire_43, N80, keyinput171);
  xnor KeyGate44 (newWire_44, N55, keyinput172);
  xor  KeyGate45 (newWire_45, N259, keyinput173);
  xor  KeyGate46 (keyNTin_Wire_1[23], N101, keyinput174);
  xnor keyNTinGate_1_23(newWire_46, keyinput271, keyNTin_Wire_1[23]);
  xor  KeyGate47 (newWire_47, N189, keyinput175);
  xor  KeyGate48 (newWire_48, N42, keyinput176);
  xnor KeyGate49 (newWire_49, N106, keyinput177);
  xor  KeyGate50 (newWire_50, N88, keyinput178);
  xor  KeyGate51 (newWire_51, N153, keyinput179);
  xor  KeyGate52 (keyNTin_Wire_1[24], N17, keyinput180);
  xor keyNTinGate_1_24(newWire_52, keyinput272, keyNTin_Wire_1[24]);
  xor  KeyGate53 (newWire_53, N146, keyinput181);
  xor  KeyGate54 (newWire_54, N87, keyinput182);
  xor  KeyGate55 (newWire_55, N51, keyinput183);
  xor  KeyGate56 (keyNTin_Wire_1[25], N29, keyinput184);
  xnor keyNTinGate_1_25(newWire_56, keyinput273, keyNTin_Wire_1[25]);
  xnor KeyGate57 (keyNTin_Wire_1[26], N255, keyinput185);
  xor keyNTinGate_1_26(KeyNOTWire_1[10], keyinput274, keyNTin_Wire_1[26]);
  not KeyNOTGate_1_10(newWire_57, KeyNOTWire_1[10]);
  xor  KeyGate58 (keyNTin_Wire_1[27], N210, keyinput186);
  xor keyNTinGate_1_27(KeyNOTWire_1[11], keyinput275, keyNTin_Wire_1[27]);
  not KeyNOTGate_1_11(newWire_58, KeyNOTWire_1[11]);
  xnor KeyGate59 (keyNTin_Wire_1[28], N171, keyinput187);
  xor keyNTinGate_1_28(KeyNOTWire_1[12], keyinput276, keyNTin_Wire_1[28]);
  not KeyNOTGate_1_12(newWire_59, KeyNOTWire_1[12]);
  xor  KeyGate60 (newWire_60, N59, keyinput188);
  xnor KeyGate61 (newWire_61, N126, keyinput189);
  xor  KeyGate62 (keyNTin_Wire_1[29], N183, keyinput190);
  xnor keyNTinGate_1_29(KeyNOTWire_1[13], keyinput277, keyNTin_Wire_1[29]);
  not KeyNOTGate_1_13(newWire_62, KeyNOTWire_1[13]);
  xnor KeyGate63 (keyNTin_Wire_1[30], N165, keyinput191);
  xor keyNTinGate_1_30(newWire_63, keyinput278, keyNTin_Wire_1[30]);
  xor  KeyGate64 (keyNTin_Wire_1[31], N156, keyinput192);
  xnor keyNTinGate_1_31(newWire_64, keyinput279, keyNTin_Wire_1[31]);
  xnor KeyGate65 (newWire_65, N237, keyinput193);
  xnor KeyGate66 (keyNTin_Wire_1[32], N8, keyinput194);
  xor keyNTinGate_1_32(KeyNOTWire_1[14], keyinput280, keyNTin_Wire_1[32]);
  not KeyNOTGate_1_14(newWire_66, KeyNOTWire_1[14]);
  xnor KeyGate67 (newWire_67, N138, keyinput195);
  xor  KeyGate68 (newWire_68, N207, keyinput196);
  xor  KeyGate69 (keyNTin_Wire_1[33], N1, keyinput197);
  xnor keyNTinGate_1_33(KeyNOTWire_1[15], keyinput281, keyNTin_Wire_1[33]);
  not KeyNOTGate_1_15(newWire_69, KeyNOTWire_1[15]);
  xnor KeyGate70 (keyNTin_Wire_1[34], N91, keyinput198);
  xor keyNTinGate_1_34(KeyNOTWire_1[16], keyinput282, keyNTin_Wire_1[34]);
  not KeyNOTGate_1_16(newWire_70, KeyNOTWire_1[16]);
  xnor KeyGate71 (newWire_71, N246, keyinput199);
  xor  KeyGate72 (newWire_72, N68, keyinput200);
  xor  KeyGate73 (keyNTin_Wire_1[35], N26, keyinput201);
  xnor keyNTinGate_1_35(newWire_73, keyinput283, keyNTin_Wire_1[35]);
  xor  KeyGate74 (newWire_74, N135, keyinput202);
  xnor KeyGate75 (newWire_75, N90, keyinput203);
  xor  KeyGate76 (newWire_76, N261, keyinput204);
  xnor KeyGate77 (newWire_77, N121, keyinput205);
  xnor KeyGate78 (keyNTin_Wire_1[36], N177, keyinput206);
  xnor keyNTinGate_1_36(KeyNOTWire_1[17], keyinput284, keyNTin_Wire_1[36]);
  not KeyNOTGate_1_17(newWire_78, KeyNOTWire_1[17]);
  xor  KeyGate79 (keyNTin_Wire_1[37], N268, keyinput207);
  xnor keyNTinGate_1_37(KeyNOTWire_1[18], keyinput285, keyNTin_Wire_1[37]);
  not KeyNOTGate_1_18(newWire_79, KeyNOTWire_1[18]);
  xor  KeyGate80 (newWire_80, N130, keyinput208);
  xor  KeyGate81 (newWire_81, N85, keyinput209);
  xnor KeyGate82 (keyNTin_Wire_1[38], N195, keyinput210);
  xnor keyNTinGate_1_38(KeyNOTWire_1[19], keyinput286, keyNTin_Wire_1[38]);
  not KeyNOTGate_1_19(newWire_82, KeyNOTWire_1[19]);
  xnor KeyGate83 (keyNTin_Wire_1[39], N36, keyinput211);
  xnor keyNTinGate_1_39(KeyNOTWire_1[20], keyinput287, keyNTin_Wire_1[39]);
  not KeyNOTGate_1_20(newWire_83, KeyNOTWire_1[20]);
  xnor KeyGate84 (keyNTin_Wire_1[40], N74, keyinput212);
  xor keyNTinGate_1_40(KeyNOTWire_1[21], keyinput288, keyNTin_Wire_1[40]);
  not KeyNOTGate_1_21(newWire_84, KeyNOTWire_1[21]);
  xor  KeyGate85 (newWire_85, N96, keyinput213);
  xnor KeyGate86 (keyNTin_Wire_1[41], N159, keyinput214);
  xnor keyNTinGate_1_41(newWire_86, keyinput289, keyNTin_Wire_1[41]);
  xor  KeyGate87 (newWire_87, N111, keyinput215);
  xnor KeyGate88 (keyNTin_Wire_1[42], N267, keyinput216);
  xor keyNTinGate_1_42(KeyNOTWire_1[22], keyinput290, keyNTin_Wire_1[42]);
  not KeyNOTGate_1_22(newWire_88, KeyNOTWire_1[22]);
  xor  KeyGate89 (keyNTin_Wire_1[43], N219, keyinput217);
  xnor keyNTinGate_1_43(newWire_89, keyinput291, keyNTin_Wire_1[43]);
  xnor KeyGate90 (keyNTin_Wire_1[44], N13, keyinput218);
  xor keyNTinGate_1_44(newWire_90, keyinput292, keyNTin_Wire_1[44]);
  xor  KeyGate91 (newWire_91, N73, keyinput219);
  xnor KeyGate92 (keyNTin_Wire_1[45], N116, keyinput220);
  xor keyNTinGate_1_45(KeyNOTWire_1[23], keyinput293, keyNTin_Wire_1[45]);
  not KeyNOTGate_1_23(newWire_92, KeyNOTWire_1[23]);
  xor  KeyGate93 (newWire_93, N143, keyinput221);
  xnor KeyGate94 (keyNTin_Wire_1[46], N260, keyinput222);
  xor keyNTinGate_1_46(newWire_94, keyinput294, keyNTin_Wire_1[46]);
  xor  KeyGate95 (newWire_95, N72, keyinput223);
  xor  KeyGate96 (keyNTin_Wire_1[47], N75, keyinput224);
  xnor keyNTinGate_1_47(newWire_96, keyinput295, keyNTin_Wire_1[47]);
  xor  KeyGate97 (newWire_97, N152, keyinput225);
  xor  KeyGate98 (newWire_98, N86, keyinput226);
  xor  KeyGate99 (newWire_99, N201, keyinput227);
  xnor KeyGate100 (newWire_100, N89, keyinput228);
  xnor KeyGate101 (keyNTin_Wire_1[48], N149, keyinput229);
  xnor keyNTinGate_1_48(newWire_101, keyinput296, keyNTin_Wire_1[48]);
  xnor KeyGate102 (newWire_102, N228, keyinput230);
  xnor KeyGate103 (newWire_103, N80, keyinput231);
  xor  KeyGate104 (keyNTin_Wire_1[49], N55, keyinput232);
  xnor keyNTinGate_1_49(newWire_104, keyinput297, keyNTin_Wire_1[49]);
  xor  KeyGate105 (keyNTin_Wire_1[50], N259, keyinput233);
  xor keyNTinGate_1_50(KeyNOTWire_1[24], keyinput298, keyNTin_Wire_1[50]);
  not KeyNOTGate_1_24(newWire_105, KeyNOTWire_1[24]);
  xor  KeyGate106 (newWire_106, N101, keyinput234);
  xnor KeyGate107 (keyNTin_Wire_1[51], N189, keyinput235);
  xnor keyNTinGate_1_51(newWire_107, keyinput299, keyNTin_Wire_1[51]);
  xor  KeyGate108 (newWire_108, N42, keyinput236);
  xor  KeyGate109 (keyNTin_Wire_1[52], N106, keyinput237);
  xor keyNTinGate_1_52(newWire_109, keyinput300, keyNTin_Wire_1[52]);
  xor  KeyGate110 (newWire_110, N88, keyinput238);
  xnor KeyGate111 (newWire_111, N153, keyinput239);
  xor  KeyGate112 (newWire_112, N17, keyinput240);
  xor  KeyGate113 (keyNTin_Wire_1[53], N146, keyinput241);
  xor keyNTinGate_1_53(newWire_113, keyinput301, keyNTin_Wire_1[53]);
  xnor KeyGate114 (keyNTin_Wire_1[54], N87, keyinput242);
  xnor keyNTinGate_1_54(newWire_114, keyinput302, keyNTin_Wire_1[54]);
  xnor KeyGate115 (keyNTin_Wire_1[55], N51, keyinput243);
  xnor keyNTinGate_1_55(newWire_115, keyinput303, keyNTin_Wire_1[55]);
  xor  KeyGate116 (newWire_116, N29, keyinput244);
  xnor KeyGate117 (keyNTin_Wire_1[56], N255, keyinput245);
  xnor keyNTinGate_1_56(newWire_117, keyinput304, keyNTin_Wire_1[56]);
  xnor KeyGate118 (newWire_118, N210, keyinput246);
  xor  KeyGate119 (keyNTin_Wire_1[57], N171, keyinput247);
  xnor keyNTinGate_1_57(KeyNOTWire_1[25], keyinput305, keyNTin_Wire_1[57]);
  not KeyNOTGate_1_25(newWire_119, KeyNOTWire_1[25]);
  and some_function (keyNTin_Wire_1[58], newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59 );
  xor keyNTinGate_1_58(newWire_120, keyinput306, keyNTin_Wire_1[58]);
  nand compl_function (keyNTin_Wire_1[59], newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83, newWire_84, newWire_85, newWire_86, newWire_87, newWire_88, newWire_89, newWire_90, newWire_91, newWire_92, newWire_93, newWire_94, newWire_95, newWire_96, newWire_97, newWire_98, newWire_99, newWire_100, newWire_101, newWire_102, newWire_103, newWire_104, newWire_105, newWire_106, newWire_107, newWire_108, newWire_109, newWire_110, newWire_111, newWire_112, newWire_113, newWire_114, newWire_115, newWire_116, newWire_117, newWire_118, newWire_119);
  xnor keyNTinGate_1_59(KeyNOTWire_1[26], keyinput307, keyNTin_Wire_1[59]);
  not KeyNOTGate_1_26(newWire_121, KeyNOTWire_1[26]);
  and finalAND (KeyWire_0_2, newWire_120, newWire_121);

endmodule /* AntiSAT */
