`timescale 1ns / 1ps
// Verilog
// c499
// Ninputs 41
// Noutputs 32
// NtotalGates 202
// XOR2 104
// AND2 40
// NOT1 40
// AND4 8
// OR4 2
// AND5 8

module top (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
                  N753,N754,N755,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
        keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
                  keyinput125, keyinput126, keyinput127,
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202,
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207,
                  keyinput208, keyinput209,
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
        keyinput250);

  input keyinput210, keyinput211, keyinput212, keyinput213, keyinput214;
  input keyinput215, keyinput216, keyinput217, keyinput218, keyinput219;
  input keyinput220, keyinput221, keyinput222, keyinput223, keyinput224;
  input keyinput225, keyinput226, keyinput227, keyinput228, keyinput229;
  input keyinput230, keyinput231, keyinput232, keyinput233, keyinput234;
  input keyinput235, keyinput236, keyinput237, keyinput238, keyinput239;
  input keyinput240, keyinput241, keyinput242, keyinput243, keyinput244;
  input keyinput245, keyinput246, keyinput247, keyinput248, keyinput249;
  input keyinput250;


  input keyinput128, keyinput129, keyinput130, keyinput131, keyinput132;
  input keyinput133, keyinput134, keyinput135, keyinput136, keyinput137;
  input keyinput138, keyinput139, keyinput140, keyinput141, keyinput142;
  input keyinput143, keyinput144, keyinput145, keyinput146, keyinput147;
  input keyinput148, keyinput149, keyinput150, keyinput151, keyinput152;
  input keyinput153, keyinput154, keyinput155, keyinput156, keyinput157;
  input keyinput158, keyinput159, keyinput160, keyinput161, keyinput162;
  input keyinput163, keyinput164, keyinput165, keyinput166, keyinput167;
  input keyinput168, keyinput169, keyinput170, keyinput171, keyinput172;
  input keyinput173, keyinput174, keyinput175, keyinput176, keyinput177;
  input keyinput178, keyinput179, keyinput180, keyinput181, keyinput182;
  input keyinput183, keyinput184, keyinput185, keyinput186, keyinput187;
  input keyinput188, keyinput189, keyinput190, keyinput191, keyinput192;
  input keyinput193, keyinput194, keyinput195, keyinput196, keyinput197;
  input keyinput198, keyinput199, keyinput200, keyinput201, keyinput202;
  input keyinput203, keyinput204, keyinput205, keyinput206, keyinput207;
  input keyinput208, keyinput209;

  wire KeyWire_0_1 , KeyWire_0_2;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31, keyinput32, keyinput33, keyinput34;
  input keyinput35, keyinput36, keyinput37, keyinput38, keyinput39;
  input keyinput40, keyinput41, keyinput42, keyinput43, keyinput44;
  input keyinput45, keyinput46, keyinput47, keyinput48, keyinput49;
  input keyinput50, keyinput51, keyinput52, keyinput53, keyinput54;
  input keyinput55, keyinput56, keyinput57, keyinput58, keyinput59;
  input keyinput60, keyinput61, keyinput62, keyinput63, keyinput64;
  input keyinput65, keyinput66, keyinput67, keyinput68, keyinput69;
  input keyinput70, keyinput71, keyinput72, keyinput73, keyinput74;
  input keyinput75, keyinput76, keyinput77, keyinput78, keyinput79;
  input keyinput80, keyinput81, keyinput82, keyinput83, keyinput84;
  input keyinput85, keyinput86, keyinput87, keyinput88, keyinput89;
  input keyinput90, keyinput91, keyinput92, keyinput93, keyinput94;
  input keyinput95, keyinput96, keyinput97, keyinput98, keyinput99;
  input keyinput100, keyinput101, keyinput102, keyinput103, keyinput104;
  input keyinput105, keyinput106, keyinput107, keyinput108, keyinput109;
  input keyinput110, keyinput111, keyinput112, keyinput113, keyinput114;
  input keyinput115, keyinput116, keyinput117, keyinput118, keyinput119;
  input keyinput120, keyinput121, keyinput122, keyinput123, keyinput124;
  input keyinput125, keyinput126, keyinput127;

  wire [0:127] keyinput_Wire_0;
  wire [0:67] KeyNOTWire_0;

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;

output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723;

  xor XOR2_1 (keyinput_Wire_0[0], N1, N5);
  xnor keyGate_0_0(KeyNOTWire_0[0], keyinput0, keyinput_Wire_0[0]);
  not KeyNOTGate_0_0(N250, KeyNOTWire_0[0]);
  xor XOR2_2 (keyinput_Wire_0[1], N9, N13);
  xnor keyGate_0_1(KeyNOTWire_0[1], keyinput1, keyinput_Wire_0[1]);
  not KeyNOTGate_0_1(N251, KeyNOTWire_0[1]);
  xor XOR2_3 (keyinput_Wire_0[2], N17, N21);
  xor keyGate_0_2(KeyNOTWire_0[2], keyinput2, keyinput_Wire_0[2]);
  not KeyNOTGate_0_2(N252, KeyNOTWire_0[2]);
  xor XOR2_4 (keyinput_Wire_0[3], N25, N29);
  xor keyGate_0_3(N253, keyinput3, keyinput_Wire_0[3]);
  xor XOR2_5 (keyinput_Wire_0[4], N33, N37);
  xnor keyGate_0_4(KeyNOTWire_0[3], keyinput4, keyinput_Wire_0[4]);
  not KeyNOTGate_0_3(N254, KeyNOTWire_0[3]);
  xor XOR2_6 (keyinput_Wire_0[5], N41, N45);
  xnor keyGate_0_5(N255, keyinput5, keyinput_Wire_0[5]);
  xor XOR2_7 (keyinput_Wire_0[6], N49, N53);
  xor keyGate_0_6(N256, keyinput6, keyinput_Wire_0[6]);
  xor XOR2_8 (keyinput_Wire_0[7], N57, N61);
  xor keyGate_0_7(N257, keyinput7, keyinput_Wire_0[7]);
  xor XOR2_9 (keyinput_Wire_0[8], N65, N69);
  xnor keyGate_0_8(N258, keyinput8, keyinput_Wire_0[8]);
  xor XOR2_10 (keyinput_Wire_0[9], N73, N77);
  xnor keyGate_0_9(KeyNOTWire_0[4], keyinput9, keyinput_Wire_0[9]);
  not KeyNOTGate_0_4(N259, KeyNOTWire_0[4]);
  xor XOR2_11 (keyinput_Wire_0[10], N81, N85);
  xnor keyGate_0_10(N260, keyinput10, keyinput_Wire_0[10]);
  xor XOR2_12 (keyinput_Wire_0[11], N89, N93);
  xor keyGate_0_11(KeyNOTWire_0[5], keyinput11, keyinput_Wire_0[11]);
  not KeyNOTGate_0_5(N261, KeyNOTWire_0[5]);
  xor XOR2_13 (keyinput_Wire_0[12], N97, N101);
  xnor keyGate_0_12(N262, keyinput12, keyinput_Wire_0[12]);
  xor XOR2_14 (keyinput_Wire_0[13], N105, N109);
  xor keyGate_0_13(KeyNOTWire_0[6], keyinput13, keyinput_Wire_0[13]);
  not KeyNOTGate_0_6(N263, KeyNOTWire_0[6]);
  xor XOR2_15 (keyinput_Wire_0[14], N113, N117);
  xor keyGate_0_14(KeyNOTWire_0[7], keyinput14, keyinput_Wire_0[14]);
  not KeyNOTGate_0_7(N264, KeyNOTWire_0[7]);
  xor XOR2_16 (keyinput_Wire_0[15], N121, N125);
  xnor keyGate_0_15(N265, keyinput15, keyinput_Wire_0[15]);
  and AND2_17 (keyinput_Wire_0[16], N129, N137);
  xnor keyGate_0_16(KeyNOTWire_0[8], keyinput16, keyinput_Wire_0[16]);
  not KeyNOTGate_0_8(N266, KeyNOTWire_0[8]);
  and AND2_18 (keyinput_Wire_0[17], N130, N137);
  xnor keyGate_0_17(KeyNOTWire_0[9], keyinput17, keyinput_Wire_0[17]);
  not KeyNOTGate_0_9(N267, KeyNOTWire_0[9]);
  and AND2_19 (keyinput_Wire_0[18], N131, N137);
  xor keyGate_0_18(KeyNOTWire_0[10], keyinput18, keyinput_Wire_0[18]);
  not KeyNOTGate_0_10(N268, KeyNOTWire_0[10]);
  and AND2_20 (keyinput_Wire_0[19], N132, N137);
  xor keyGate_0_19(KeyNOTWire_0[11], keyinput19, keyinput_Wire_0[19]);
  not KeyNOTGate_0_11(N269, KeyNOTWire_0[11]);
  and AND2_21 (keyinput_Wire_0[20], N133, N137);
  xor keyGate_0_20(KeyNOTWire_0[12], keyinput20, keyinput_Wire_0[20]);
  not KeyNOTGate_0_12(N270, KeyNOTWire_0[12]);
  and AND2_22 (keyinput_Wire_0[21], N134, N137);
  xor keyGate_0_21(KeyNOTWire_0[13], keyinput21, keyinput_Wire_0[21]);
  not KeyNOTGate_0_13(N271, KeyNOTWire_0[13]);
  and AND2_23 (keyinput_Wire_0[22], N135, N137);
  xnor keyGate_0_22(KeyNOTWire_0[14], keyinput22, keyinput_Wire_0[22]);
  not KeyNOTGate_0_14(N272, KeyNOTWire_0[14]);
  and AND2_24 (keyinput_Wire_0[23], N136, N137);
  xnor keyGate_0_23(KeyNOTWire_0[15], keyinput23, keyinput_Wire_0[23]);
  not KeyNOTGate_0_15(N273, KeyNOTWire_0[15]);
  xor XOR2_25 (keyinput_Wire_0[24], N1, N17);
  xnor keyGate_0_24(N274, keyinput24, keyinput_Wire_0[24]);
  xor XOR2_26 (keyinput_Wire_0[25], N33, N49);
  xnor keyGate_0_25(N275, keyinput25, keyinput_Wire_0[25]);
  xor XOR2_27 (keyinput_Wire_0[26], N5, N21);
  xnor keyGate_0_26(N276, keyinput26, keyinput_Wire_0[26]);
  xor XOR2_28 (keyinput_Wire_0[27], N37, N53);
  xor keyGate_0_27(KeyNOTWire_0[16], keyinput27, keyinput_Wire_0[27]);
  not KeyNOTGate_0_16(N277, KeyNOTWire_0[16]);
  xor XOR2_29 (keyinput_Wire_0[28], N9, N25);
  xnor keyGate_0_28(N278, keyinput28, keyinput_Wire_0[28]);
  xor XOR2_30 (keyinput_Wire_0[29], N41, N57);
  xor keyGate_0_29(KeyNOTWire_0[17], keyinput29, keyinput_Wire_0[29]);
  not KeyNOTGate_0_17(N279, KeyNOTWire_0[17]);
  xor XOR2_31 (keyinput_Wire_0[30], N13, N29);
  xor keyGate_0_30(KeyNOTWire_0[18], keyinput30, keyinput_Wire_0[30]);
  not KeyNOTGate_0_18(N280, KeyNOTWire_0[18]);
  xor XOR2_32 (keyinput_Wire_0[31], N45, N61);
  xor keyGate_0_31(KeyNOTWire_0[19], keyinput31, keyinput_Wire_0[31]);
  not KeyNOTGate_0_19(N281, KeyNOTWire_0[19]);
  xor XOR2_33 (keyinput_Wire_0[32], N65, N81);
  xor keyGate_0_32(N282, keyinput32, keyinput_Wire_0[32]);
  xor XOR2_34 (keyinput_Wire_0[33], N97, N113);
  xor keyGate_0_33(N283, keyinput33, keyinput_Wire_0[33]);
  xor XOR2_35 (keyinput_Wire_0[34], N69, N85);
  xor keyGate_0_34(N284, keyinput34, keyinput_Wire_0[34]);
  xor XOR2_36 (keyinput_Wire_0[35], N101, N117);
  xor keyGate_0_35(KeyNOTWire_0[20], keyinput35, keyinput_Wire_0[35]);
  not KeyNOTGate_0_20(N285, KeyNOTWire_0[20]);
  xor XOR2_37 (keyinput_Wire_0[36], N73, N89);
  xnor keyGate_0_36(KeyNOTWire_0[21], keyinput36, keyinput_Wire_0[36]);
  not KeyNOTGate_0_21(N286, KeyNOTWire_0[21]);
  xor XOR2_38 (keyinput_Wire_0[37], N105, N121);
  xnor keyGate_0_37(N287, keyinput37, keyinput_Wire_0[37]);
  xor XOR2_39 (keyinput_Wire_0[38], N77, N93);
  xor keyGate_0_38(N288, keyinput38, keyinput_Wire_0[38]);
  xor XOR2_40 (keyinput_Wire_0[39], N109, N125);
  xor keyGate_0_39(N289, keyinput39, keyinput_Wire_0[39]);
  xor XOR2_41 (keyinput_Wire_0[40], N250, N251);
  xnor keyGate_0_40(N290, keyinput40, keyinput_Wire_0[40]);
  xor XOR2_42 (keyinput_Wire_0[41], N252, N253);
  xor keyGate_0_41(KeyNOTWire_0[22], keyinput41, keyinput_Wire_0[41]);
  not KeyNOTGate_0_22(N293, KeyNOTWire_0[22]);
  xor XOR2_43 (keyinput_Wire_0[42], N254, N255);
  xnor keyGate_0_42(KeyNOTWire_0[23], keyinput42, keyinput_Wire_0[42]);
  not KeyNOTGate_0_23(N296, KeyNOTWire_0[23]);
  xor XOR2_44 (keyinput_Wire_0[43], N256, N257);
  xor keyGate_0_43(N299, keyinput43, keyinput_Wire_0[43]);
  xor XOR2_45 (keyinput_Wire_0[44], N258, N259);
  xor keyGate_0_44(N302, keyinput44, keyinput_Wire_0[44]);
  xor XOR2_46 (keyinput_Wire_0[45], N260, N261);
  xnor keyGate_0_45(N305, keyinput45, keyinput_Wire_0[45]);
  xor XOR2_47 (keyinput_Wire_0[46], N262, N263);
  xor keyGate_0_46(N308, keyinput46, keyinput_Wire_0[46]);
  xor XOR2_48 (keyinput_Wire_0[47], N264, N265);
  xor keyGate_0_47(KeyNOTWire_0[24], keyinput47, keyinput_Wire_0[47]);
  not KeyNOTGate_0_24(N311, KeyNOTWire_0[24]);
  xor XOR2_49 (keyinput_Wire_0[48], N274, N275);
  xnor keyGate_0_48(KeyNOTWire_0[25], keyinput48, keyinput_Wire_0[48]);
  not KeyNOTGate_0_25(N314, KeyNOTWire_0[25]);
  xor XOR2_50 (keyinput_Wire_0[49], N276, N277);
  xor keyGate_0_49(N315, keyinput49, keyinput_Wire_0[49]);
  xor XOR2_51 (keyinput_Wire_0[50], N278, N279);
  xnor keyGate_0_50(N316, keyinput50, keyinput_Wire_0[50]);
  xor XOR2_52 (keyinput_Wire_0[51], N280, N281);
  xor keyGate_0_51(KeyNOTWire_0[26], keyinput51, keyinput_Wire_0[51]);
  not KeyNOTGate_0_26(N317, KeyNOTWire_0[26]);
  xor XOR2_53 (keyinput_Wire_0[52], N282, N283);
  xnor keyGate_0_52(N318, keyinput52, keyinput_Wire_0[52]);
  xor XOR2_54 (keyinput_Wire_0[53], N284, N285);
  xnor keyGate_0_53(N319, keyinput53, keyinput_Wire_0[53]);
  xor XOR2_55 (keyinput_Wire_0[54], N286, N287);
  xnor keyGate_0_54(N320, keyinput54, keyinput_Wire_0[54]);
  xor XOR2_56 (keyinput_Wire_0[55], N288, N289);
  xor keyGate_0_55(KeyNOTWire_0[27], keyinput55, keyinput_Wire_0[55]);
  not KeyNOTGate_0_27(N321, KeyNOTWire_0[27]);
  xor XOR2_57 (keyinput_Wire_0[56], N290, N293);
  xor keyGate_0_56(KeyNOTWire_0[28], keyinput56, keyinput_Wire_0[56]);
  not KeyNOTGate_0_28(N338, KeyNOTWire_0[28]);
  xor XOR2_58 (keyinput_Wire_0[57], N296, N299);
  xor keyGate_0_57(N339, keyinput57, keyinput_Wire_0[57]);
  xor XOR2_59 (keyinput_Wire_0[58], N290, N296);
  xnor keyGate_0_58(KeyNOTWire_0[29], keyinput58, keyinput_Wire_0[58]);
  not KeyNOTGate_0_29(N340, KeyNOTWire_0[29]);
  xor XOR2_60 (keyinput_Wire_0[59], N293, N299);
  xor keyGate_0_59(N341, keyinput59, keyinput_Wire_0[59]);
  xor XOR2_61 (keyinput_Wire_0[60], N302, N305);
  xnor keyGate_0_60(KeyNOTWire_0[30], keyinput60, keyinput_Wire_0[60]);
  not KeyNOTGate_0_30(N342, KeyNOTWire_0[30]);
  xor XOR2_62 (keyinput_Wire_0[61], N308, N311);
  xnor keyGate_0_61(N343, keyinput61, keyinput_Wire_0[61]);
  xor XOR2_63 (keyinput_Wire_0[62], N302, N308);
  xnor keyGate_0_62(N344, keyinput62, keyinput_Wire_0[62]);
  xor XOR2_64 (keyinput_Wire_0[63], N305, N311);
  xor keyGate_0_63(KeyNOTWire_0[31], keyinput63, keyinput_Wire_0[63]);
  not KeyNOTGate_0_31(N345, KeyNOTWire_0[31]);
  xor XOR2_65 (keyinput_Wire_0[64], N266, N342);
  xnor keyGate_0_64(KeyNOTWire_0[32], keyinput64, keyinput_Wire_0[64]);
  not KeyNOTGate_0_32(N346, KeyNOTWire_0[32]);
  xor XOR2_66 (keyinput_Wire_0[65], N267, N343);
  xor keyGate_0_65(N347, keyinput65, keyinput_Wire_0[65]);
  xor XOR2_67 (keyinput_Wire_0[66], N268, N344);
  xor keyGate_0_66(N348, keyinput66, keyinput_Wire_0[66]);
  xor XOR2_68 (keyinput_Wire_0[67], N269, N345);
  xnor keyGate_0_67(N349, keyinput67, keyinput_Wire_0[67]);
  xor XOR2_69 (keyinput_Wire_0[68], N270, N338);
  xnor keyGate_0_68(N350, keyinput68, keyinput_Wire_0[68]);
  xor XOR2_70 (keyinput_Wire_0[69], N271, N339);
  xnor keyGate_0_69(KeyNOTWire_0[33], keyinput69, keyinput_Wire_0[69]);
  not KeyNOTGate_0_33(N351, KeyNOTWire_0[33]);
  xor XOR2_71 (keyinput_Wire_0[70], N272, N340);
  xnor keyGate_0_70(KeyNOTWire_0[34], keyinput70, keyinput_Wire_0[70]);
  not KeyNOTGate_0_34(N352, KeyNOTWire_0[34]);
  xor XOR2_72 (keyinput_Wire_0[71], N273, N341);
  xnor keyGate_0_71(KeyNOTWire_0[35], keyinput71, keyinput_Wire_0[71]);
  not KeyNOTGate_0_35(N353, KeyNOTWire_0[35]);
  xor XOR2_73 (keyinput_Wire_0[72], N314, N346);
  xor keyGate_0_72(KeyNOTWire_0[36], keyinput72, keyinput_Wire_0[72]);
  not KeyNOTGate_0_36(N354, KeyNOTWire_0[36]);
  xor XOR2_74 (keyinput_Wire_0[73], N315, N347);
  xnor keyGate_0_73(N367, keyinput73, keyinput_Wire_0[73]);
  xor XOR2_75 (keyinput_Wire_0[74], N316, N348);
  xor keyGate_0_74(KeyNOTWire_0[37], keyinput74, keyinput_Wire_0[74]);
  not KeyNOTGate_0_37(N380, KeyNOTWire_0[37]);
  xor XOR2_76 (keyinput_Wire_0[75], N317, N349);
  xnor keyGate_0_75(KeyNOTWire_0[38], keyinput75, keyinput_Wire_0[75]);
  not KeyNOTGate_0_38(N393, KeyNOTWire_0[38]);
  xor XOR2_77 (keyinput_Wire_0[76], N318, N350);
  xnor keyGate_0_76(KeyNOTWire_0[39], keyinput76, keyinput_Wire_0[76]);
  not KeyNOTGate_0_39(N406, KeyNOTWire_0[39]);
  xor XOR2_78 (keyinput_Wire_0[77], N319, N351);
  xnor keyGate_0_77(KeyNOTWire_0[40], keyinput77, keyinput_Wire_0[77]);
  not KeyNOTGate_0_40(N419, KeyNOTWire_0[40]);
  xor XOR2_79 (keyinput_Wire_0[78], N320, N352);
  xnor keyGate_0_78(N432, keyinput78, keyinput_Wire_0[78]);
  xor XOR2_80 (keyinput_Wire_0[79], N321, N353);
  xor keyGate_0_79(KeyNOTWire_0[41], keyinput79, keyinput_Wire_0[79]);
  not KeyNOTGate_0_41(N445, KeyNOTWire_0[41]);
  not NOT1_81 (keyinput_Wire_0[80], N354);
  xor keyGate_0_80(KeyNOTWire_0[42], keyinput80, keyinput_Wire_0[80]);
  not KeyNOTGate_0_42(N554, KeyNOTWire_0[42]);
not NOT1_82 (N555, N367);
not NOT1_83 (N556, N380);
not NOT1_84 (N557, N354);
not NOT1_85 (N558, N367);
  not NOT1_86 (keyinput_Wire_0[81], N393);
  xor keyGate_0_81(KeyNOTWire_0[43], keyinput81, keyinput_Wire_0[81]);
  not KeyNOTGate_0_43(N559, KeyNOTWire_0[43]);
not NOT1_87 (N560, N354);
not NOT1_88 (N561, N380);
not NOT1_89 (N562, N393);
not NOT1_90 (N563, N367);
not NOT1_91 (N564, N380);
not NOT1_92 (N565, N393);
not NOT1_93 (N566, N419);
not NOT1_94 (N567, N445);
not NOT1_95 (N568, N419);
not NOT1_96 (N569, N432);
not NOT1_97 (N570, N406);
not NOT1_98 (N571, N445);
not NOT1_99 (N572, N406);
not NOT1_100 (N573, N432);
  not NOT1_101 (keyinput_Wire_0[82], N406);
  xor keyGate_0_82(N574, keyinput82, keyinput_Wire_0[82]);
  not NOT1_102 (keyinput_Wire_0[83], N419);
  xor keyGate_0_83(N575, keyinput83, keyinput_Wire_0[83]);
  not NOT1_103 (keyinput_Wire_0[84], N432);
  xnor keyGate_0_84(N576, keyinput84, keyinput_Wire_0[84]);
  not NOT1_104 (keyinput_Wire_0[85], N406);
  xor keyGate_0_85(N577, keyinput85, keyinput_Wire_0[85]);
  not NOT1_105 (keyinput_Wire_0[86], N419);
  xnor keyGate_0_86(KeyNOTWire_0[44], keyinput86, keyinput_Wire_0[86]);
  not KeyNOTGate_0_44(N578, KeyNOTWire_0[44]);
  not NOT1_106 (keyinput_Wire_0[87], N445);
  xor keyGate_0_87(KeyNOTWire_0[45], keyinput87, keyinput_Wire_0[87]);
  not KeyNOTGate_0_45(N579, KeyNOTWire_0[45]);
  not NOT1_107 (keyinput_Wire_0[88], N406);
  xor keyGate_0_88(KeyNOTWire_0[46], keyinput88, keyinput_Wire_0[88]);
  not KeyNOTGate_0_46(N580, KeyNOTWire_0[46]);
  not NOT1_108 (keyinput_Wire_0[89], N432);
  xnor keyGate_0_89(N581, keyinput89, keyinput_Wire_0[89]);
  not NOT1_109 (keyinput_Wire_0[90], N445);
  xor keyGate_0_90(N582, keyinput90, keyinput_Wire_0[90]);
  not NOT1_110 (keyinput_Wire_0[91], N419);
  xnor keyGate_0_91(KeyNOTWire_0[47], keyinput91, keyinput_Wire_0[91]);
  not KeyNOTGate_0_47(N583, KeyNOTWire_0[47]);
  not NOT1_111 (keyinput_Wire_0[92], N432);
  xnor keyGate_0_92(KeyNOTWire_0[48], keyinput92, keyinput_Wire_0[92]);
  not KeyNOTGate_0_48(N584, KeyNOTWire_0[48]);
  not NOT1_112 (keyinput_Wire_0[93], N445);
  xor keyGate_0_93(N585, keyinput93, keyinput_Wire_0[93]);
not NOT1_113 (N586, N367);
  not NOT1_114 (keyinput_Wire_0[94], N393);
  xor keyGate_0_94(N587, keyinput94, keyinput_Wire_0[94]);
not NOT1_115 (N588, N367);
not NOT1_116 (N589, N380);
not NOT1_117 (N590, N354);
not NOT1_118 (N591, N393);
not NOT1_119 (N592, N354);
not NOT1_120 (N593, N380);
  and AND4_121 (keyinput_Wire_0[95], N554, N555, N556, N393);
  xor keyGate_0_95(N594, keyinput95, keyinput_Wire_0[95]);
and AND4_122 (N595, N557, N558, N380, N559);
and AND4_123 (N596, N560, N367, N561, N562);
and AND4_124 (N597, N354, N563, N564, N565);
  and AND4_125 (keyinput_Wire_0[96], N574, N575, N576, N445);
  xor keyGate_0_96(KeyNOTWire_0[49], keyinput96, keyinput_Wire_0[96]);
  not KeyNOTGate_0_49(N598, KeyNOTWire_0[49]);
  and AND4_126 (keyinput_Wire_0[97], N577, N578, N432, N579);
  xor keyGate_0_97(N599, keyinput97, keyinput_Wire_0[97]);
  and AND4_127 (keyinput_Wire_0[98], N580, N419, N581, N582);
  xnor keyGate_0_98(KeyNOTWire_0[50], keyinput98, keyinput_Wire_0[98]);
  not KeyNOTGate_0_50(N600, KeyNOTWire_0[50]);
  and AND4_128 (keyinput_Wire_0[99], N406, N583, N584, N585);
  xnor keyGate_0_99(KeyNOTWire_0[51], keyinput99, keyinput_Wire_0[99]);
  not KeyNOTGate_0_51(N601, KeyNOTWire_0[51]);
or OR4_129 (N602, N594, N595, N596, N597);
  or OR4_130 (keyinput_Wire_0[100], N598, N599, N600, N601);
  xnor keyGate_0_100(N607, keyinput100, keyinput_Wire_0[100]);
and AND5_131 (N620, N406, N566, N432, N567, N602);
  and AND5_132 (keyinput_Wire_0[101], N406, N568, N569, N445, N602);
  xnor keyGate_0_101(N625, keyinput101, keyinput_Wire_0[101]);
  and AND5_133 (keyinput_Wire_0[102], N570, N419, N432, N571, N602);
  xor keyGate_0_102(KeyNOTWire_0[52], keyinput102, keyinput_Wire_0[102]);
  not KeyNOTGate_0_52(N630, KeyNOTWire_0[52]);
and AND5_134 (N635, N572, N419, N573, N445, N602);
and AND5_135 (N640, N354, N586, N380, N587, N607);
and AND5_136 (N645, N354, N588, N589, N393, N607);
and AND5_137 (N650, N590, N367, N380, N591, N607);
and AND5_138 (N655, N592, N367, N593, N393, N607);
and AND2_139 (N692, N354, N620);
and AND2_140 (N693, N367, N620);
and AND2_141 (N694, N380, N620);
and AND2_142 (N695, N393, N620);
and AND2_143 (N696, N354, N625);
and AND2_144 (N697, N367, N625);
and AND2_145 (N698, N380, N625);
and AND2_146 (N699, N393, N625);
and AND2_147 (N700, N354, N630);
and AND2_148 (N701, N367, N630);
and AND2_149 (N702, N380, N630);
and AND2_150 (N703, N393, N630);
and AND2_151 (N704, N354, N635);
and AND2_152 (N705, N367, N635);
and AND2_153 (N706, N380, N635);
and AND2_154 (N707, N393, N635);
and AND2_155 (N708, N406, N640);
  and AND2_156 (keyinput_Wire_0[103], N419, N640);
  xor keyGate_0_103(KeyNOTWire_0[53], keyinput103, keyinput_Wire_0[103]);
  not KeyNOTGate_0_53(N709, KeyNOTWire_0[53]);
and AND2_157 (N710, N432, N640);
and AND2_158 (N711, N445, N640);
  and AND2_159 (keyinput_Wire_0[104], N406, N645);
  xnor keyGate_0_104(KeyNOTWire_0[54], keyinput104, keyinput_Wire_0[104]);
  not KeyNOTGate_0_54(N712, KeyNOTWire_0[54]);
and AND2_160 (N713, N419, N645);
and AND2_161 (N714, N432, N645);
and AND2_162 (N715, N445, N645);
and AND2_163 (N716, N406, N650);
and AND2_164 (N717, N419, N650);
and AND2_165 (N718, N432, N650);
and AND2_166 (N719, N445, N650);
and AND2_167 (N720, N406, N655);
and AND2_168 (N721, N419, N655);
and AND2_169 (N722, N432, N655);
and AND2_170 (N723, N445, N655);
  xor XOR2_171 (keyinput_Wire_0[105], N1, N692);
  xor keyGate_0_105(N724, keyinput105, keyinput_Wire_0[105]);
xor XOR2_172 (N725, N5, N693);
  xor XOR2_173 (keyinput_Wire_0[106], N9, N694);
  xnor keyGate_0_106(N726, keyinput106, keyinput_Wire_0[106]);
xor XOR2_174 (N727, N13, N695);
  xor XOR2_175 (keyinput_Wire_0[107], N17, N696);
  xor keyGate_0_107(KeyNOTWire_0[55], keyinput107, keyinput_Wire_0[107]);
  not KeyNOTGate_0_55(KeyWire_0_1, KeyNOTWire_0[55]);
  xor flip_it (N728, KeyWire_0_1, KeyWire_0_2 );
  xor XOR2_176 (keyinput_Wire_0[108], N21, N697);
  xnor keyGate_0_108(KeyNOTWire_0[56], keyinput108, keyinput_Wire_0[108]);
  not KeyNOTGate_0_56(N729, KeyNOTWire_0[56]);
  xor XOR2_177 (keyinput_Wire_0[109], N25, N698);
  xnor keyGate_0_109(KeyNOTWire_0[57], keyinput109, keyinput_Wire_0[109]);
  not KeyNOTGate_0_57(N730, KeyNOTWire_0[57]);
  xor XOR2_178 (keyinput_Wire_0[110], N29, N699);
  xor keyGate_0_110(N731, keyinput110, keyinput_Wire_0[110]);
  xor XOR2_179 (keyinput_Wire_0[111], N33, N700);
  xor keyGate_0_111(KeyNOTWire_0[58], keyinput111, keyinput_Wire_0[111]);
  not KeyNOTGate_0_58(N732, KeyNOTWire_0[58]);
  xor XOR2_180 (keyinput_Wire_0[112], N37, N701);
  xor keyGate_0_112(N733, keyinput112, keyinput_Wire_0[112]);
  xor XOR2_181 (keyinput_Wire_0[113], N41, N702);
  xnor keyGate_0_113(KeyNOTWire_0[59], keyinput113, keyinput_Wire_0[113]);
  not KeyNOTGate_0_59(N734, KeyNOTWire_0[59]);
  xor XOR2_182 (keyinput_Wire_0[114], N45, N703);
  xor keyGate_0_114(KeyNOTWire_0[60], keyinput114, keyinput_Wire_0[114]);
  not KeyNOTGate_0_60(N735, KeyNOTWire_0[60]);
  xor XOR2_183 (keyinput_Wire_0[115], N49, N704);
  xnor keyGate_0_115(N736, keyinput115, keyinput_Wire_0[115]);
xor XOR2_184 (N737, N53, N705);
  xor XOR2_185 (keyinput_Wire_0[116], N57, N706);
  xnor keyGate_0_116(KeyNOTWire_0[61], keyinput116, keyinput_Wire_0[116]);
  not KeyNOTGate_0_61(N738, KeyNOTWire_0[61]);
  xor XOR2_186 (keyinput_Wire_0[117], N61, N707);
  xor keyGate_0_117(KeyNOTWire_0[62], keyinput117, keyinput_Wire_0[117]);
  not KeyNOTGate_0_62(N739, KeyNOTWire_0[62]);
  xor XOR2_187 (keyinput_Wire_0[118], N65, N708);
  xnor keyGate_0_118(N740, keyinput118, keyinput_Wire_0[118]);
  xor XOR2_188 (keyinput_Wire_0[119], N69, N709);
  xor keyGate_0_119(N741, keyinput119, keyinput_Wire_0[119]);
  xor XOR2_189 (keyinput_Wire_0[120], N73, N710);
  xnor keyGate_0_120(KeyNOTWire_0[63], keyinput120, keyinput_Wire_0[120]);
  not KeyNOTGate_0_63(N742, KeyNOTWire_0[63]);
xor XOR2_190 (N743, N77, N711);
  xor XOR2_191 (keyinput_Wire_0[121], N81, N712);
  xnor keyGate_0_121(KeyNOTWire_0[64], keyinput121, keyinput_Wire_0[121]);
  not KeyNOTGate_0_64(N744, KeyNOTWire_0[64]);
xor XOR2_192 (N745, N85, N713);
xor XOR2_193 (N746, N89, N714);
  xor XOR2_194 (keyinput_Wire_0[122], N93, N715);
  xor keyGate_0_122(KeyNOTWire_0[65], keyinput122, keyinput_Wire_0[122]);
  not KeyNOTGate_0_65(N747, KeyNOTWire_0[65]);
  xor XOR2_195 (keyinput_Wire_0[123], N97, N716);
  xnor keyGate_0_123(N748, keyinput123, keyinput_Wire_0[123]);
  xor XOR2_196 (keyinput_Wire_0[124], N101, N717);
  xnor keyGate_0_124(N749, keyinput124, keyinput_Wire_0[124]);
xor XOR2_197 (N750, N105, N718);
  xor XOR2_198 (keyinput_Wire_0[125], N109, N719);
  xor keyGate_0_125(KeyNOTWire_0[66], keyinput125, keyinput_Wire_0[125]);
  not KeyNOTGate_0_66(N751, KeyNOTWire_0[66]);
  xor XOR2_199 (keyinput_Wire_0[126], N113, N720);
  xnor keyGate_0_126(N752, keyinput126, keyinput_Wire_0[126]);
  xor XOR2_200 (keyinput_Wire_0[127], N117, N721);
  xnor keyGate_0_127(KeyNOTWire_0[67], keyinput127, keyinput_Wire_0[127]);
  not KeyNOTGate_0_67(N753, KeyNOTWire_0[67]);
xor XOR2_201 (N754, N121, N722);
xor XOR2_202 (N755, N125, N723);

AntiSAT some_name( KeyWire_0_2, N25, N5, N136, N93, N109, N132, N135, N37, N137, N125, N117, N53, N45, N65, N9, N49, N29, N69, N33, N121, N131, N130, N17, N41, N73, N13, N134, N97, N113, N1, N129, N105, N101, N61, N85, N89, N133, N81, N57, N21, N77, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
       keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
       keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
       keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
       keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
       keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
       keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
       keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
       keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
       keyinput250);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N25, N5, N136, N93, N109, N132, N135, N37, N137, N125, N117, N53, N45, N65, N9, N49, N29, N69, N33, N121, N131, N130, N17, N41, N73, N13, N134, N97, N113, N1, N129, N105, N101, N61, N85, N89, N133, N81, N57, N21, N77, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, keyinput208, keyinput209 ,
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
        keyinput250);

  input keyinput210, keyinput211, keyinput212, keyinput213, keyinput214;
  input keyinput215, keyinput216, keyinput217, keyinput218, keyinput219;
  input keyinput220, keyinput221, keyinput222, keyinput223, keyinput224;
  input keyinput225, keyinput226, keyinput227, keyinput228, keyinput229;
  input keyinput230, keyinput231, keyinput232, keyinput233, keyinput234;
  input keyinput235, keyinput236, keyinput237, keyinput238, keyinput239;
  input keyinput240, keyinput241, keyinput242, keyinput243, keyinput244;
  input keyinput245, keyinput246, keyinput247, keyinput248, keyinput249;
  input keyinput250;

  wire [0:40] keyNTin_Wire_1;
  wire [0:20] KeyNOTWire_1;

  input N25, N5, N136, N93, N109, N132, N135, N37, N137, N125, N117, N53, N45, N65, N9, N49, N29, N69, N33, N121, N131, N130, N17, N41, N73, N13, N134, N97, N113, N1, N129, N105, N101, N61, N85, N89, N133, N81, N57, N21, N77;
  input keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, keyinput208, keyinput209;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83 ;

  xor  KeyGate0 (newWire_0, N25, keyinput128);
  xnor KeyGate1 (newWire_1, N5, keyinput129);
  xnor KeyGate2 (keyNTin_Wire_1[0], N136, keyinput130);
  xor keyNTinGate_1_0(newWire_2, keyinput210, keyNTin_Wire_1[0]);
  xnor KeyGate3 (keyNTin_Wire_1[1], N93, keyinput131);
  xnor keyNTinGate_1_1(newWire_3, keyinput211, keyNTin_Wire_1[1]);
  xor  KeyGate4 (keyNTin_Wire_1[2], N109, keyinput132);
  xor keyNTinGate_1_2(KeyNOTWire_1[0], keyinput212, keyNTin_Wire_1[2]);
  not KeyNOTGate_1_0(newWire_4, KeyNOTWire_1[0]);
  xor  KeyGate5 (newWire_5, N132, keyinput133);
  xnor KeyGate6 (newWire_6, N135, keyinput134);
  xnor KeyGate7 (keyNTin_Wire_1[3], N37, keyinput135);
  xnor keyNTinGate_1_3(newWire_7, keyinput213, keyNTin_Wire_1[3]);
  xnor KeyGate8 (newWire_8, N137, keyinput136);
  xnor KeyGate9 (keyNTin_Wire_1[4], N125, keyinput137);
  xnor keyNTinGate_1_4(newWire_9, keyinput214, keyNTin_Wire_1[4]);
  xor  KeyGate10 (keyNTin_Wire_1[5], N117, keyinput138);
  xor keyNTinGate_1_5(KeyNOTWire_1[1], keyinput215, keyNTin_Wire_1[5]);
  not KeyNOTGate_1_1(newWire_10, KeyNOTWire_1[1]);
  xnor KeyGate11 (newWire_11, N53, keyinput139);
  xor  KeyGate12 (keyNTin_Wire_1[6], N45, keyinput140);
  xor keyNTinGate_1_6(KeyNOTWire_1[2], keyinput216, keyNTin_Wire_1[6]);
  not KeyNOTGate_1_2(newWire_12, KeyNOTWire_1[2]);
  xor  KeyGate13 (newWire_13, N65, keyinput141);
  xor  KeyGate14 (keyNTin_Wire_1[7], N9, keyinput142);
  xor keyNTinGate_1_7(KeyNOTWire_1[3], keyinput217, keyNTin_Wire_1[7]);
  not KeyNOTGate_1_3(newWire_14, KeyNOTWire_1[3]);
  xnor KeyGate15 (keyNTin_Wire_1[8], N49, keyinput143);
  xnor keyNTinGate_1_8(KeyNOTWire_1[4], keyinput218, keyNTin_Wire_1[8]);
  not KeyNOTGate_1_4(newWire_15, KeyNOTWire_1[4]);
  xor  KeyGate16 (keyNTin_Wire_1[9], N29, keyinput144);
  xor keyNTinGate_1_9(KeyNOTWire_1[5], keyinput219, keyNTin_Wire_1[9]);
  not KeyNOTGate_1_5(newWire_16, KeyNOTWire_1[5]);
  xnor KeyGate17 (keyNTin_Wire_1[10], N69, keyinput145);
  xnor keyNTinGate_1_10(newWire_17, keyinput220, keyNTin_Wire_1[10]);
  xnor KeyGate18 (newWire_18, N33, keyinput146);
  xnor KeyGate19 (keyNTin_Wire_1[11], N121, keyinput147);
  xnor keyNTinGate_1_11(KeyNOTWire_1[6], keyinput221, keyNTin_Wire_1[11]);
  not KeyNOTGate_1_6(newWire_19, KeyNOTWire_1[6]);
  xor  KeyGate20 (keyNTin_Wire_1[12], N131, keyinput148);
  xor keyNTinGate_1_12(KeyNOTWire_1[7], keyinput222, keyNTin_Wire_1[12]);
  not KeyNOTGate_1_7(newWire_20, KeyNOTWire_1[7]);
  xnor KeyGate21 (newWire_21, N130, keyinput149);
  xnor KeyGate22 (keyNTin_Wire_1[13], N17, keyinput150);
  xnor keyNTinGate_1_13(newWire_22, keyinput223, keyNTin_Wire_1[13]);
  xnor KeyGate23 (newWire_23, N41, keyinput151);
  xor  KeyGate24 (newWire_24, N73, keyinput152);
  xor  KeyGate25 (keyNTin_Wire_1[14], N13, keyinput153);
  xor keyNTinGate_1_14(newWire_25, keyinput224, keyNTin_Wire_1[14]);
  xor  KeyGate26 (keyNTin_Wire_1[15], N134, keyinput154);
  xor keyNTinGate_1_15(newWire_26, keyinput225, keyNTin_Wire_1[15]);
  xor  KeyGate27 (newWire_27, N97, keyinput155);
  xor  KeyGate28 (newWire_28, N113, keyinput156);
  xor  KeyGate29 (keyNTin_Wire_1[16], N1, keyinput157);
  xnor keyNTinGate_1_16(newWire_29, keyinput226, keyNTin_Wire_1[16]);
  xnor KeyGate30 (newWire_30, N129, keyinput158);
  xor  KeyGate31 (keyNTin_Wire_1[17], N105, keyinput159);
  xnor keyNTinGate_1_17(newWire_31, keyinput227, keyNTin_Wire_1[17]);
  xor  KeyGate32 (newWire_32, N101, keyinput160);
  xnor KeyGate33 (keyNTin_Wire_1[18], N61, keyinput161);
  xnor keyNTinGate_1_18(KeyNOTWire_1[8], keyinput228, keyNTin_Wire_1[18]);
  not KeyNOTGate_1_8(newWire_33, KeyNOTWire_1[8]);
  xor  KeyGate34 (keyNTin_Wire_1[19], N85, keyinput162);
  xor keyNTinGate_1_19(newWire_34, keyinput229, keyNTin_Wire_1[19]);
  xor  KeyGate35 (newWire_35, N89, keyinput163);
  xor  KeyGate36 (keyNTin_Wire_1[20], N133, keyinput164);
  xnor keyNTinGate_1_20(KeyNOTWire_1[9], keyinput230, keyNTin_Wire_1[20]);
  not KeyNOTGate_1_9(newWire_36, KeyNOTWire_1[9]);
  xnor KeyGate37 (keyNTin_Wire_1[21], N81, keyinput165);
  xor keyNTinGate_1_21(KeyNOTWire_1[10], keyinput231, keyNTin_Wire_1[21]);
  not KeyNOTGate_1_10(newWire_37, KeyNOTWire_1[10]);
  xor  KeyGate38 (keyNTin_Wire_1[22], N57, keyinput166);
  xnor keyNTinGate_1_22(KeyNOTWire_1[11], keyinput232, keyNTin_Wire_1[22]);
  not KeyNOTGate_1_11(newWire_38, KeyNOTWire_1[11]);
  xor  KeyGate39 (newWire_39, N21, keyinput167);
  xor  KeyGate40 (newWire_40, N77, keyinput168);
  xor  KeyGate41 (newWire_41, N25, keyinput169);
  xor  KeyGate42 (newWire_42, N5, keyinput170);
  xor  KeyGate43 (keyNTin_Wire_1[23], N136, keyinput171);
  xor keyNTinGate_1_23(KeyNOTWire_1[12], keyinput233, keyNTin_Wire_1[23]);
  not KeyNOTGate_1_12(newWire_43, KeyNOTWire_1[12]);
  xor  KeyGate44 (newWire_44, N93, keyinput172);
  xor  KeyGate45 (keyNTin_Wire_1[24], N109, keyinput173);
  xnor keyNTinGate_1_24(newWire_45, keyinput234, keyNTin_Wire_1[24]);
  xnor KeyGate46 (newWire_46, N132, keyinput174);
  xnor KeyGate47 (newWire_47, N135, keyinput175);
  xor  KeyGate48 (newWire_48, N37, keyinput176);
  xnor KeyGate49 (keyNTin_Wire_1[25], N137, keyinput177);
  xor keyNTinGate_1_25(KeyNOTWire_1[13], keyinput235, keyNTin_Wire_1[25]);
  not KeyNOTGate_1_13(newWire_49, KeyNOTWire_1[13]);
  xnor KeyGate50 (newWire_50, N125, keyinput178);
  xnor KeyGate51 (keyNTin_Wire_1[26], N117, keyinput179);
  xnor keyNTinGate_1_26(newWire_51, keyinput236, keyNTin_Wire_1[26]);
  xnor KeyGate52 (keyNTin_Wire_1[27], N53, keyinput180);
  xor keyNTinGate_1_27(KeyNOTWire_1[14], keyinput237, keyNTin_Wire_1[27]);
  not KeyNOTGate_1_14(newWire_52, KeyNOTWire_1[14]);
  xnor KeyGate53 (keyNTin_Wire_1[28], N45, keyinput181);
  xor keyNTinGate_1_28(KeyNOTWire_1[15], keyinput238, keyNTin_Wire_1[28]);
  not KeyNOTGate_1_15(newWire_53, KeyNOTWire_1[15]);
  xnor KeyGate54 (newWire_54, N65, keyinput182);
  xor  KeyGate55 (keyNTin_Wire_1[29], N9, keyinput183);
  xor keyNTinGate_1_29(newWire_55, keyinput239, keyNTin_Wire_1[29]);
  xnor KeyGate56 (newWire_56, N49, keyinput184);
  xor  KeyGate57 (newWire_57, N29, keyinput185);
  xnor KeyGate58 (newWire_58, N69, keyinput186);
  xnor KeyGate59 (newWire_59, N33, keyinput187);
  xnor KeyGate60 (newWire_60, N121, keyinput188);
  xor  KeyGate61 (newWire_61, N131, keyinput189);
  xor  KeyGate62 (newWire_62, N130, keyinput190);
  xnor KeyGate63 (keyNTin_Wire_1[30], N17, keyinput191);
  xor keyNTinGate_1_30(KeyNOTWire_1[16], keyinput240, keyNTin_Wire_1[30]);
  not KeyNOTGate_1_16(newWire_63, KeyNOTWire_1[16]);
  xor  KeyGate64 (newWire_64, N41, keyinput192);
  xnor KeyGate65 (keyNTin_Wire_1[31], N73, keyinput193);
  xnor keyNTinGate_1_31(newWire_65, keyinput241, keyNTin_Wire_1[31]);
  xnor KeyGate66 (keyNTin_Wire_1[32], N13, keyinput194);
  xor keyNTinGate_1_32(KeyNOTWire_1[17], keyinput242, keyNTin_Wire_1[32]);
  not KeyNOTGate_1_17(newWire_66, KeyNOTWire_1[17]);
  xor  KeyGate67 (keyNTin_Wire_1[33], N134, keyinput195);
  xnor keyNTinGate_1_33(KeyNOTWire_1[18], keyinput243, keyNTin_Wire_1[33]);
  not KeyNOTGate_1_18(newWire_67, KeyNOTWire_1[18]);
  xnor KeyGate68 (keyNTin_Wire_1[34], N97, keyinput196);
  xor keyNTinGate_1_34(newWire_68, keyinput244, keyNTin_Wire_1[34]);
  xor  KeyGate69 (newWire_69, N113, keyinput197);
  xnor KeyGate70 (newWire_70, N1, keyinput198);
  xor  KeyGate71 (newWire_71, N129, keyinput199);
  xnor KeyGate72 (keyNTin_Wire_1[35], N105, keyinput200);
  xnor keyNTinGate_1_35(KeyNOTWire_1[19], keyinput245, keyNTin_Wire_1[35]);
  not KeyNOTGate_1_19(newWire_72, KeyNOTWire_1[19]);
  xnor KeyGate73 (keyNTin_Wire_1[36], N101, keyinput201);
  xnor keyNTinGate_1_36(newWire_73, keyinput246, keyNTin_Wire_1[36]);
  xor  KeyGate74 (newWire_74, N61, keyinput202);
  xor  KeyGate75 (keyNTin_Wire_1[37], N85, keyinput203);
  xnor keyNTinGate_1_37(newWire_75, keyinput247, keyNTin_Wire_1[37]);
  xnor KeyGate76 (newWire_76, N89, keyinput204);
  xnor KeyGate77 (newWire_77, N133, keyinput205);
  xnor KeyGate78 (newWire_78, N81, keyinput206);
  xnor KeyGate79 (newWire_79, N57, keyinput207);
  xor  KeyGate80 (keyNTin_Wire_1[38], N21, keyinput208);
  xor keyNTinGate_1_38(newWire_80, keyinput248, keyNTin_Wire_1[38]);
  xor  KeyGate81 (newWire_81, N77, keyinput209);
  and some_function (newWire_82, newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40 );
  nand compl_function (keyNTin_Wire_1[39], newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81);
  xor keyNTinGate_1_39(newWire_83, keyinput249, keyNTin_Wire_1[39]);
  and finalAND (keyNTin_Wire_1[40], newWire_82, newWire_83);
  xor keyNTinGate_1_40(KeyNOTWire_1[20], keyinput250, keyNTin_Wire_1[40]);
  not KeyNOTGate_1_20(KeyWire_0_2, KeyNOTWire_1[20]);

endmodule /* AntiSAT */
