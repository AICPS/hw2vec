// Verilog File 
module top (G1gat,G8gat,G13gat,G17gat,G26gat,G29gat,G36gat,G42gat,G51gat,
G55gat,G59gat,G68gat,G72gat,G73gat,G74gat,G75gat,G80gat,G85gat,G86gat,
G87gat,G88gat,G89gat,G90gat,G91gat,G96gat,G101gat,G106gat,G111gat,G116gat,
G121gat,G126gat,G130gat,G135gat,G138gat,G143gat,G146gat,G149gat,G152gat,G153gat,
G156gat,G159gat,G165gat,G171gat,G177gat,G183gat,G189gat,G195gat,G201gat,G207gat,
G210gat,G219gat,G228gat,G237gat,G246gat,G255gat,G259gat,G260gat,G261gat,G267gat,
G268gat,G388gat,G389gat,G390gat,G391gat,G418gat,G419gat,G420gat,G421gat,G422gat,
G423gat,G446gat,G447gat,G448gat,G449gat,G450gat,G767gat,G768gat,G850gat,G863gat,
G864gat,G865gat,G866gat,G874gat,G878gat,G879gat,G880gat,keyinput0,keyinput1,keyinput2,
keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,
keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,
keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,
keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,
keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,
keyinput53,keyinput54,keyinput55,keyinput56,keyinput57,keyinput58);

input G1gat,G8gat,G13gat,G17gat,G26gat,G29gat,G36gat,G42gat,G51gat,
G55gat,G59gat,G68gat,G72gat,G73gat,G74gat,G75gat,G80gat,G85gat,G86gat,
G87gat,G88gat,G89gat,G90gat,G91gat,G96gat,G101gat,G106gat,G111gat,G116gat,
G121gat,G126gat,G130gat,G135gat,G138gat,G143gat,G146gat,G149gat,G152gat,G153gat,
G156gat,G159gat,G165gat,G171gat,G177gat,G183gat,G189gat,G195gat,G201gat,G207gat,
G210gat,G219gat,G228gat,G237gat,G246gat,G255gat,G259gat,G260gat,G261gat,G267gat,
G268gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,
keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,
keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,
keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,keyinput38,
keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,keyinput48,
keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,keyinput55,keyinput56,keyinput57,keyinput58;

output G388gat,G389gat,G390gat,G391gat,G418gat,G419gat,G420gat,G421gat,G422gat,
G423gat,G446gat,G447gat,G448gat,G449gat,G450gat,G767gat,G768gat,G850gat,G863gat,
G864gat,G865gat,G866gat,G874gat,G878gat,G879gat,G880gat;

wire G269gat,G270gat,G273gat,G276gat,G279gat,G280gat,G284gat,G285gat,G286gat,
G287gat,G290gat,G291gat,G292gat,G293gat,G294gat,G295gat,G296gat,G297gat,G298gat,
G301gat,G302gat,G303gat,G304gat,G305gat,G306gat,G307gat,G308gat,G309gat,G310gat,
G316gat,G317gat,G318gat,G319gat,G322gat,G323gat,G324gat,G325gat,G326gat,G327gat,
G328gat,G329gat,G330gat,G331gat,G332gat,G333gat,G334gat,G335gat,G336gat,G337gat,
G338gat,G339gat,G340gat,G341gat,G342gat,G343gat,G344gat,G345gat,G346gat,G347gat,
G348gat,G349gat,G350gat,G351gat,G352gat,G353gat,G354gat,G355gat,G356gat,G357gat,
G360gat,G363gat,G366gat,G369gat,G375gat,G376gat,G379gat,G382gat,G385gat,G392gat,
G393gat,G399gat,G400gat,G401gat,G402gat,G403gat,G404gat,G405gat,G406gat,G407gat,
G408gat,G409gat,G410gat,G411gat,G412gat,G413gat,G414gat,G415gat,G416gat,G417gat,
G424gat,G425gat,G426gat,G427gat,G432gat,G437gat,G442gat,G443gat,G444gat,G445gat,
G451gat,G460gat,G463gat,G466gat,G475gat,G476gat,G477gat,G478gat,G479gat,G480gat,
G481gat,G482gat,G483gat,G488gat,G489gat,G490gat,G491gat,G492gat,G495gat,G498gat,
G499gat,G500gat,G501gat,G502gat,G503gat,G504gat,G505gat,G506gat,G507gat,G508gat,
G509gat,G510gat,G511gat,G512gat,G513gat,G514gat,G515gat,G516gat,G517gat,G518gat,
G519gat,G520gat,G521gat,G522gat,G523gat,G524gat,G525gat,G526gat,G527gat,G528gat,
G529gat,G530gat,G533gat,G536gat,G537gat,G538gat,G539gat,G540gat,G541gat,G542gat,
G543gat,G544gat,G547gat,G550gat,G551gat,G552gat,G553gat,G557gat,G561gat,G565gat,
G569gat,G573gat,G577gat,G581gat,G585gat,G586gat,G587gat,G588gat,G589gat,G590gat,
G593gat,G596gat,G597gat,G600gat,G605gat,G606gat,G609gat,G615gat,G616gat,G619gat,
G624gat,G625gat,G628gat,G631gat,G632gat,G635gat,G640gat,G641gat,G644gat,G650gat,
G651gat,G654gat,G659gat,G660gat,G661gat,G662gat,G665gat,G669gat,G670gat,G673gat,
G677gat,G678gat,G682gat,G686gat,G687gat,G692gat,G696gat,G697gat,G700gat,G704gat,
G705gat,G708gat,G712gat,G713gat,G717gat,G721gat,G722gat,G727gat,G731gat,G732gat,
G733gat,G734gat,G735gat,G736gat,G737gat,G738gat,G739gat,G740gat,G741gat,G742gat,
G743gat,G744gat,G745gat,G746gat,G747gat,G748gat,G749gat,G750gat,G751gat,G752gat,
G753gat,G754gat,G755gat,G756gat,G757gat,G758gat,G759gat,G760gat,G761gat,G762gat,
G763gat,G764gat,G765gat,G766gat,G769gat,G770gat,G771gat,G772gat,G773gat,G777gat,
G778gat,G781gat,G782gat,G785gat,G786gat,G787gat,G788gat,G789gat,G790gat,G791gat,
G792gat,G793gat,G794gat,G795gat,G796gat,G802gat,G803gat,G804gat,G805gat,G806gat,
G807gat,G808gat,G809gat,G810gat,G811gat,G812gat,G813gat,G814gat,G815gat,G819gat,
G822gat,G825gat,G826gat,G827gat,G828gat,G829gat,G830gat,G831gat,G832gat,G833gat,
G834gat,G835gat,G836gat,G837gat,G838gat,G839gat,G840gat,G841gat,G842gat,G843gat,
G844gat,G845gat,G846gat,G847gat,G848gat,G849gat,G851gat,G852gat,G853gat,G854gat,
G855gat,G856gat,G857gat,G858gat,G859gat,G860gat,G861gat,G862gat,G867gat,G868gat,
G869gat,G870gat,G871gat,G872gat,G873gat,G875gat,G876gat,G877gat,muxed0,muxed1,
muxed2,muxed3,muxed4,muxed5,muxed6,muxed7,muxed8,muxed9,muxed10,muxed11,
muxed12,muxed13,muxed14,muxed15,muxed16,muxed17,muxed18,muxed19,muxed20,muxed21,
muxed22,muxed23,muxed24,muxed25,muxed26,muxed27,muxed28,muxed29,muxed30,muxed31,
muxed32,muxed33,muxed34,muxed35,muxed36,muxed37,muxed38,muxed39,muxed40,muxed41,
muxed42,muxed43,muxed44,muxed45,muxed46,muxed47,muxed48,muxed49,muxed50,muxed51,
muxed52,muxed53,muxed54,muxed55,muxed56,muxed57,muxed58;
nand gate_0(G269gat,G1gat,G8gat,G13gat,G17gat);
nand gate_1(G270gat,G1gat,G26gat,G13gat,G17gat);
and gate_2(G273gat,G29gat,G36gat,G42gat);
and gate_3(G276gat,G1gat,G26gat,G51gat);
nand gate_4(G279gat,G1gat,G8gat,G51gat,G17gat);
nand gate_5(G280gat,G1gat,G8gat,G13gat,G55gat);
nand gate_6(G284gat,G59gat,G42gat,G68gat,G72gat);
nand gate_7(G285gat,G29gat,G68gat);
nand gate_8(G286gat,G59gat,G68gat,G74gat);
and gate_9(G287gat,G29gat,G75gat,G80gat);
and gate_10(G290gat,G29gat,G75gat,G42gat);
and gate_11(G291gat,G29gat,G36gat,G80gat);
and gate_12(G292gat,G29gat,G36gat,G42gat);
and gate_13(G293gat,G59gat,G75gat,G80gat);
and gate_14(G294gat,G59gat,G75gat,G42gat);
and gate_15(G295gat,G59gat,G36gat,G80gat);
and gate_16(G296gat,G59gat,G36gat,G42gat);
and gate_17(G297gat,G85gat,G86gat);
or gate_18(G298gat,G87gat,G88gat);
nand gate_19(G301gat,G91gat,G96gat);
or gate_20(G302gat,G91gat,G96gat);
nand gate_21(G303gat,G101gat,G106gat);
or gate_22(G304gat,G101gat,G106gat);
nand gate_23(G305gat,G111gat,G116gat);
or gate_24(G306gat,G111gat,G116gat);
nand gate_25(G307gat,G121gat,G126gat);
or gate_26(G308gat,G121gat,G126gat);
and gate_27(G309gat,G8gat,G138gat);
not gate_28(G310gat,G268gat);
and gate_29(G316gat,G51gat,G138gat);
and gate_30(G317gat,G17gat,G138gat);
and gate_31(G318gat,G152gat,G138gat);
nand gate_32(G319gat,G59gat,G156gat);
nor gate_33(G322gat,G17gat,G42gat);
and gate_34(G323gat,G17gat,G42gat);
nand gate_35(G324gat,G159gat,G165gat);
or gate_36(G325gat,G159gat,G165gat);
nand gate_37(G326gat,G171gat,G177gat);
or gate_38(G327gat,G171gat,G177gat);
nand gate_39(G328gat,G183gat,G189gat);
or gate_40(G329gat,G183gat,G189gat);
nand gate_41(G330gat,G195gat,G201gat);
or gate_42(G331gat,G195gat,G201gat);
and gate_43(G332gat,G210gat,G91gat);
and gate_44(G333gat,G210gat,G96gat);
and gate_45(G334gat,G210gat,G101gat);
and gate_46(G335gat,G210gat,G106gat);
and gate_47(G336gat,G210gat,G111gat);
and gate_48(G337gat,G255gat,G259gat);
and gate_49(G338gat,G210gat,G116gat);
and gate_50(G339gat,G255gat,G260gat);
and gate_51(G340gat,G210gat,G121gat);
and gate_52(G341gat,G255gat,G267gat);
not gate_53(G342gat,G269gat);
not gate_54(G343gat,G273gat);
or gate_55(G344gat,G270gat,G273gat);
not gate_56(G345gat,G276gat);
not gate_57(G346gat,G276gat);
not gate_58(G347gat,muxed53);
nor gate_59(G348gat,G280gat,muxed46);
or gate_60(G349gat,G280gat,G285gat);
or gate_61(G350gat,G280gat,G286gat);
not gate_62(G351gat,G293gat);
not gate_63(G352gat,G294gat);
not gate_64(G353gat,G295gat);
not gate_65(G354gat,G296gat);
nand gate_66(G355gat,G89gat,muxed4);
and gate_67(G356gat,G90gat,muxed4);
nand gate_68(G357gat,muxed16,G302gat);
nand gate_69(G360gat,muxed0,G304gat);
nand gate_70(G363gat,G305gat,G306gat);
nand gate_71(G366gat,muxed6,G308gat);
not gate_72(G369gat,G310gat);
nor gate_73(G375gat,G322gat,G323gat);
nand gate_74(G376gat,G324gat,G325gat);
nand gate_75(G379gat,G326gat,G327gat);
nand gate_76(G382gat,G328gat,G329gat);
nand gate_77(G385gat,G330gat,G331gat);
buf gate_78(G388gat,G290gat);
buf gate_79(G389gat,G291gat);
buf gate_80(G390gat,G292gat);
buf gate_81(G391gat,G297gat);
or gate_82(G392gat,G270gat,G343gat);
not gate_83(G393gat,G345gat);
not gate_84(G399gat,G346gat);
and gate_85(G400gat,G348gat,G73gat);
not gate_86(G401gat,G349gat);
not gate_87(G402gat,G350gat);
not gate_88(G403gat,G355gat);
not gate_89(G404gat,G357gat);
not gate_90(G405gat,muxed13);
and gate_91(G406gat,G357gat,muxed13);
not gate_92(G407gat,G363gat);
not gate_93(G408gat,G366gat);
and gate_94(G409gat,G363gat,G366gat);
nand gate_95(G410gat,G347gat,G352gat);
not gate_96(G411gat,muxed44);
not gate_97(G412gat,G379gat);
and gate_98(G413gat,muxed44,G379gat);
not gate_99(G414gat,G382gat);
not gate_100(G415gat,G385gat);
and gate_101(G416gat,G382gat,G385gat);
and gate_102(G417gat,G210gat,G369gat);
buf gate_103(G418gat,G342gat);
buf gate_104(G419gat,G344gat);
buf gate_105(G420gat,G351gat);
buf gate_106(G421gat,G353gat);
buf gate_107(G422gat,muxed9);
buf gate_108(G423gat,G356gat);
not gate_109(G424gat,G400gat);
and gate_110(G425gat,G404gat,G405gat);
and gate_111(G426gat,G407gat,G408gat);
and gate_112(G427gat,G319gat,G393gat,G55gat);
and gate_113(G432gat,G393gat,G17gat,G287gat);
nand gate_114(G437gat,G393gat,G287gat,G55gat);
nand gate_115(G442gat,G375gat,G59gat,G156gat,G393gat);
nand gate_116(G443gat,G393gat,G319gat,G17gat);
and gate_117(G444gat,muxed57,G412gat);
and gate_118(G445gat,G414gat,G415gat);
buf gate_119(G446gat,G392gat);
buf gate_120(G447gat,G399gat);
buf gate_121(G448gat,G401gat);
buf gate_122(G449gat,G402gat);
buf gate_123(G450gat,G403gat);
not gate_124(G451gat,G424gat);
nor gate_125(G460gat,muxed11,G425gat);
nor gate_126(G463gat,G409gat,G426gat);
nand gate_127(G466gat,G442gat,G410gat);
and gate_128(G475gat,G143gat,G427gat);
and gate_129(G476gat,G310gat,G432gat);
and gate_130(G477gat,G146gat,G427gat);
and gate_131(G478gat,G310gat,G432gat);
and gate_132(G479gat,G149gat,G427gat);
and gate_133(G480gat,G310gat,G432gat);
and gate_134(G481gat,G153gat,G427gat);
and gate_135(G482gat,G310gat,G432gat);
nand gate_136(G483gat,G443gat,G1gat);
or gate_137(G488gat,G369gat,G437gat);
or gate_138(G489gat,G369gat,G437gat);
or gate_139(G490gat,G369gat,G437gat);
or gate_140(G491gat,G369gat,G437gat);
nor gate_141(G492gat,G413gat,muxed55);
nor gate_142(G495gat,G416gat,G445gat);
nand gate_143(G498gat,G130gat,muxed10);
or gate_144(G499gat,G130gat,muxed10);
nand gate_145(G500gat,G463gat,G135gat);
or gate_146(G501gat,G463gat,G135gat);
and gate_147(G502gat,G91gat,G466gat);
nor gate_148(G503gat,G475gat,G476gat);
and gate_149(G504gat,G96gat,G466gat);
nor gate_150(G505gat,G477gat,G478gat);
and gate_151(G506gat,G101gat,G466gat);
nor gate_152(G507gat,G479gat,G480gat);
and gate_153(G508gat,G106gat,G466gat);
nor gate_154(G509gat,G481gat,G482gat);
and gate_155(G510gat,G143gat,G483gat);
and gate_156(G511gat,G111gat,G466gat);
and gate_157(G512gat,G146gat,G483gat);
and gate_158(G513gat,G116gat,G466gat);
and gate_159(G514gat,G149gat,G483gat);
and gate_160(G515gat,G121gat,G466gat);
and gate_161(G516gat,G153gat,G483gat);
and gate_162(G517gat,G126gat,G466gat);
nand gate_163(G518gat,G130gat,muxed54);
or gate_164(G519gat,G130gat,muxed54);
nand gate_165(G520gat,G495gat,G207gat);
or gate_166(G521gat,G495gat,G207gat);
and gate_167(G522gat,G451gat,G159gat);
and gate_168(G523gat,G451gat,G165gat);
and gate_169(G524gat,G451gat,G171gat);
and gate_170(G525gat,G451gat,G177gat);
and gate_171(G526gat,G451gat,G183gat);
nand gate_172(G527gat,G451gat,G189gat);
nand gate_173(G528gat,G451gat,G195gat);
nand gate_174(G529gat,G451gat,G201gat);
nand gate_175(G530gat,G498gat,muxed8);
nand gate_176(G533gat,muxed41,G501gat);
nor gate_177(G536gat,G309gat,G502gat);
nor gate_178(G537gat,G316gat,G504gat);
nor gate_179(G538gat,G317gat,G506gat);
nor gate_180(G539gat,G318gat,G508gat);
nor gate_181(G540gat,G510gat,G511gat);
nor gate_182(G541gat,G512gat,G513gat);
nor gate_183(G542gat,G514gat,G515gat);
nor gate_184(G543gat,G516gat,G517gat);
nand gate_185(G544gat,G518gat,muxed52);
nand gate_186(G547gat,G520gat,G521gat);
not gate_187(G550gat,muxed7);
not gate_188(G551gat,G533gat);
and gate_189(G552gat,muxed7,G533gat);
nand gate_190(G553gat,G536gat,G503gat);
nand gate_191(G557gat,G537gat,G505gat);
nand gate_192(G561gat,G538gat,G507gat);
nand gate_193(G565gat,G539gat,G509gat);
nand gate_194(G569gat,G488gat,G540gat);
nand gate_195(G573gat,G489gat,G541gat);
nand gate_196(G577gat,G490gat,muxed38);
nand gate_197(G581gat,G491gat,G543gat);
not gate_198(G585gat,muxed51);
not gate_199(G586gat,G547gat);
and gate_200(G587gat,muxed51,G547gat);
and gate_201(G588gat,G550gat,G551gat);
and gate_202(G589gat,G585gat,G586gat);
nand gate_203(G590gat,G553gat,G159gat);
or gate_204(G593gat,G553gat,G159gat);
and gate_205(G596gat,G246gat,G553gat);
nand gate_206(G597gat,G557gat,G165gat);
or gate_207(G600gat,G557gat,G165gat);
and gate_208(G605gat,G246gat,G557gat);
nand gate_209(G606gat,G561gat,G171gat);
or gate_210(G609gat,G561gat,G171gat);
and gate_211(G615gat,G246gat,G561gat);
nand gate_212(G616gat,G565gat,G177gat);
or gate_213(G619gat,G565gat,G177gat);
and gate_214(G624gat,G246gat,G565gat);
nand gate_215(G625gat,G569gat,G183gat);
or gate_216(G628gat,G569gat,G183gat);
and gate_217(G631gat,G246gat,G569gat);
nand gate_218(G632gat,G573gat,G189gat);
or gate_219(G635gat,G573gat,G189gat);
and gate_220(G640gat,G246gat,G573gat);
nand gate_221(G641gat,G577gat,G195gat);
or gate_222(G644gat,G577gat,G195gat);
and gate_223(G650gat,G246gat,G577gat);
nand gate_224(G651gat,G581gat,G201gat);
or gate_225(G654gat,G581gat,G201gat);
and gate_226(G659gat,G246gat,G581gat);
nor gate_227(G660gat,muxed5,G588gat);
nor gate_228(G661gat,muxed49,G589gat);
not gate_229(G662gat,muxed12);
and gate_230(G665gat,G593gat,muxed12);
nor gate_231(G669gat,G596gat,muxed36);
not gate_232(G670gat,G597gat);
and gate_233(G673gat,G600gat,G597gat);
nor gate_234(G677gat,G605gat,G523gat);
not gate_235(G678gat,G606gat);
and gate_236(G682gat,G609gat,G606gat);
nor gate_237(G686gat,G615gat,G524gat);
not gate_238(G687gat,G616gat);
and gate_239(G692gat,G619gat,G616gat);
nor gate_240(G696gat,G624gat,G525gat);
not gate_241(G697gat,G625gat);
and gate_242(G700gat,G628gat,G625gat);
nor gate_243(G704gat,G631gat,G526gat);
not gate_244(G705gat,G632gat);
and gate_245(G708gat,muxed31,G632gat);
nor gate_246(G712gat,G337gat,G640gat);
not gate_247(G713gat,G641gat);
and gate_248(G717gat,G644gat,G641gat);
nor gate_249(G721gat,G339gat,G650gat);
not gate_250(G722gat,G651gat);
and gate_251(G727gat,G654gat,G651gat);
nor gate_252(G731gat,G341gat,G659gat);
nand gate_253(G732gat,G654gat,G261gat);
nand gate_254(G733gat,G644gat,G654gat,G261gat);
nand gate_255(G734gat,muxed31,G644gat,G654gat,G261gat);
not gate_256(G735gat,G662gat);
and gate_257(G736gat,G228gat,G665gat);
and gate_258(G737gat,G237gat,G662gat);
not gate_259(G738gat,G670gat);
and gate_260(G739gat,G228gat,G673gat);
and gate_261(G740gat,G237gat,G670gat);
not gate_262(G741gat,G678gat);
and gate_263(G742gat,G228gat,G682gat);
and gate_264(G743gat,G237gat,G678gat);
not gate_265(G744gat,G687gat);
and gate_266(G745gat,G228gat,muxed14);
and gate_267(G746gat,G237gat,G687gat);
not gate_268(G747gat,G697gat);
and gate_269(G748gat,G228gat,G700gat);
and gate_270(G749gat,G237gat,G697gat);
not gate_271(G750gat,G705gat);
and gate_272(G751gat,G228gat,muxed43);
and gate_273(G752gat,G237gat,G705gat);
not gate_274(G753gat,G713gat);
and gate_275(G754gat,G228gat,G717gat);
and gate_276(G755gat,G237gat,G713gat);
not gate_277(G756gat,G722gat);
nor gate_278(G757gat,G727gat,G261gat);
and gate_279(G758gat,G727gat,G261gat);
and gate_280(G759gat,G228gat,G727gat);
and gate_281(G760gat,G237gat,G722gat);
nand gate_282(G761gat,G644gat,G722gat);
nand gate_283(G762gat,muxed31,G713gat);
nand gate_284(G763gat,muxed31,G644gat,G722gat);
nand gate_285(G764gat,G609gat,G687gat);
nand gate_286(G765gat,G600gat,G678gat);
nand gate_287(G766gat,G600gat,G609gat,G687gat);
buf gate_288(G767gat,muxed3);
buf gate_289(G768gat,muxed47);
nor gate_290(G769gat,G736gat,G737gat);
nor gate_291(G770gat,G739gat,G740gat);
nor gate_292(G771gat,G742gat,G743gat);
nor gate_293(G772gat,G745gat,G746gat);
nand gate_294(G773gat,muxed50,G762gat,G763gat,G734gat);
nor gate_295(G777gat,G748gat,G749gat);
nand gate_296(G778gat,G753gat,G761gat,G733gat);
nor gate_297(G781gat,G751gat,G752gat);
nand gate_298(G782gat,G756gat,G732gat);
nor gate_299(G785gat,G754gat,G755gat);
nor gate_300(G786gat,muxed18,G758gat);
nor gate_301(G787gat,G759gat,G760gat);
nor gate_302(G788gat,G700gat,G773gat);
and gate_303(G789gat,G700gat,G773gat);
nor gate_304(G790gat,muxed43,muxed22);
and gate_305(G791gat,muxed43,muxed22);
nor gate_306(G792gat,G717gat,G782gat);
and gate_307(G793gat,G717gat,G782gat);
and gate_308(G794gat,G219gat,G786gat);
nand gate_309(G795gat,G628gat,G773gat);
nand gate_310(G796gat,G795gat,G747gat);
nor gate_311(G802gat,G788gat,G789gat);
nor gate_312(G803gat,G790gat,muxed42);
nor gate_313(G804gat,G792gat,G793gat);
nor gate_314(G805gat,G340gat,G794gat);
nor gate_315(G806gat,muxed14,G796gat);
and gate_316(G807gat,muxed14,G796gat);
and gate_317(G808gat,G219gat,G802gat);
and gate_318(G809gat,G219gat,G803gat);
and gate_319(G810gat,G219gat,G804gat);
nand gate_320(G811gat,G805gat,G787gat,G731gat,G529gat);
nand gate_321(G812gat,G619gat,G796gat);
nand gate_322(G813gat,G609gat,G619gat,G796gat);
nand gate_323(G814gat,G600gat,G609gat,G619gat,G796gat);
nand gate_324(G815gat,G738gat,G765gat,G766gat,G814gat);
nand gate_325(G819gat,G741gat,G764gat,G813gat);
nand gate_326(G822gat,G744gat,muxed26);
nor gate_327(G825gat,muxed29,G807gat);
nor gate_328(G826gat,G335gat,G808gat);
nor gate_329(G827gat,G336gat,G809gat);
nor gate_330(G828gat,G338gat,G810gat);
not gate_331(G829gat,G811gat);
nor gate_332(G830gat,G665gat,G815gat);
and gate_333(G831gat,G665gat,G815gat);
nor gate_334(G832gat,G673gat,G819gat);
and gate_335(G833gat,G673gat,G819gat);
nor gate_336(G834gat,G682gat,G822gat);
and gate_337(G835gat,G682gat,G822gat);
and gate_338(G836gat,G219gat,muxed27);
nand gate_339(G837gat,G826gat,G777gat,G704gat);
nand gate_340(G838gat,muxed34,G781gat,G712gat,G527gat);
nand gate_341(G839gat,G828gat,G785gat,G721gat,G528gat);
not gate_342(G840gat,G829gat);
nand gate_343(G841gat,G815gat,G593gat);
nor gate_344(G842gat,G830gat,G831gat);
nor gate_345(G843gat,G832gat,muxed20);
nor gate_346(G844gat,G834gat,G835gat);
nor gate_347(G845gat,G334gat,muxed40);
not gate_348(G846gat,muxed48);
not gate_349(G847gat,muxed30);
not gate_350(G848gat,G839gat);
and gate_351(G849gat,G735gat,G841gat);
buf gate_352(G850gat,G840gat);
and gate_353(G851gat,G219gat,muxed37);
and gate_354(G852gat,G219gat,G843gat);
and gate_355(G853gat,G219gat,G844gat);
nand gate_356(G854gat,muxed23,G772gat,G696gat);
not gate_357(G855gat,G846gat);
not gate_358(G856gat,G847gat);
not gate_359(G857gat,G848gat);
not gate_360(G858gat,G849gat);
nor gate_361(G859gat,G417gat,muxed35);
nor gate_362(G860gat,G332gat,G852gat);
nor gate_363(G861gat,muxed28,G853gat);
not gate_364(G862gat,muxed21);
buf gate_365(G863gat,G855gat);
buf gate_366(G864gat,G856gat);
buf gate_367(G865gat,G857gat);
buf gate_368(G866gat,G858gat);
nand gate_369(G867gat,muxed33,G769gat,G669gat);
nand gate_370(G868gat,G860gat,muxed56,G677gat);
nand gate_371(G869gat,G861gat,G771gat,G686gat);
not gate_372(G870gat,muxed19);
not gate_373(G871gat,muxed32);
not gate_374(G872gat,G868gat);
not gate_375(G873gat,G869gat);
buf gate_376(G874gat,muxed17);
not gate_377(G875gat,G871gat);
not gate_378(G876gat,G872gat);
not gate_379(G877gat,G873gat);
buf gate_380(G878gat,G875gat);
buf gate_381(G879gat,G876gat);
buf gate_382(G880gat,muxed2);
assign muxed0 = keyinput0 ? G303gat : muxed1;
assign muxed1 = keyinput1 ? G767gat : G297gat;
assign muxed2 = keyinput2 ? G877gat : G767gat;
assign muxed3 = keyinput3 ? G660gat : G306gat;
assign muxed4 = keyinput4 ? G298gat : G660gat;
assign muxed5 = keyinput5 ? G552gat : muxed41;
assign muxed6 = keyinput6 ? G307gat : G552gat;
assign muxed7 = keyinput7 ? G530gat : G803gat;
assign muxed8 = keyinput8 ? G499gat : G758gat;
assign muxed9 = keyinput9 ? G354gat : G499gat;
assign muxed10 = keyinput10 ? G460gat : G414gat;
assign muxed11 = keyinput11 ? G406gat : G366gat;
assign muxed12 = keyinput12 ? G590gat : G406gat;
assign muxed13 = keyinput13 ? G360gat : G871gat;
assign muxed14 = keyinput14 ? G692gat : muxed15;
assign muxed15 = keyinput15 ? G874gat : G692gat;
assign muxed16 = keyinput16 ? G301gat : G874gat;
assign muxed17 = keyinput17 ? G870gat : G766gat;
assign muxed18 = keyinput18 ? G757gat : G870gat;
assign muxed19 = keyinput19 ? G862gat : G835gat;
assign muxed20 = keyinput20 ? G833gat : G862gat;
assign muxed21 = keyinput21 ? G854gat : G855gat;
assign muxed22 = keyinput22 ? G778gat : G854gat;
assign muxed23 = keyinput23 ? muxed39 : G445gat;
assign muxed24 = keyinput24 ? G842gat : muxed39;
assign muxed25 = keyinput25 ? G836gat : muxed42;
assign muxed26 = keyinput26 ? G812gat : G836gat;
assign muxed27 = keyinput27 ? G825gat : G463gat;
assign muxed28 = keyinput28 ? G333gat : G825gat;
assign muxed29 = keyinput29 ? G806gat : G406gat;
assign muxed30 = keyinput30 ? G838gat : G806gat;
assign muxed31 = keyinput31 ? G635gat : muxed32;
assign muxed32 = keyinput32 ? G867gat : G831gat;
assign muxed33 = keyinput33 ? G859gat : G734gat;
assign muxed34 = keyinput34 ? G827gat : G859gat;
assign muxed35 = keyinput35 ? G851gat : G297gat;
assign muxed36 = keyinput36 ? G522gat : G851gat;
assign muxed37 = keyinput37 ? muxed24 : G836gat;
assign muxed38 = keyinput38 ? G542gat : muxed24;
assign muxed39 = keyinput39 ? G845gat : G834gat;
assign muxed40 = keyinput40 ? muxed25 : G862gat;
assign muxed41 = keyinput41 ? G500gat : muxed25;
assign muxed42 = keyinput42 ? G791gat : G751gat;
assign muxed43 = keyinput43 ? G708gat : G392gat;
assign muxed44 = keyinput44 ? G376gat : muxed45;
assign muxed45 = keyinput45 ? G768gat : G735gat;
assign muxed46 = keyinput46 ? G284gat : G768gat;
assign muxed47 = keyinput47 ? G661gat : G552gat;
assign muxed48 = keyinput48 ? G837gat : G661gat;
assign muxed49 = keyinput49 ? muxed58 : G778gat;
assign muxed50 = keyinput50 ? G750gat : muxed58;
assign muxed51 = keyinput51 ? G544gat : G869gat;
assign muxed52 = keyinput52 ? G519gat : G867gat;
assign muxed53 = keyinput53 ? G279gat : G519gat;
assign muxed54 = keyinput54 ? G492gat : G596gat;
assign muxed55 = keyinput55 ? G444gat : G852gat;
assign muxed56 = keyinput56 ? G770gat : G444gat;
assign muxed57 = keyinput57 ? G411gat : G721gat;
assign muxed58 = keyinput58 ? G587gat : G411gat;
endmodule
