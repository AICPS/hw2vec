`timescale 1ns / 1ps
// Verilog
// c432
// Ninputs 36
// Noutputs 7
// NtotalGates 160
// NOT1 40
// NAND2 64
// NOR2 19
// AND9 3
// XOR2 18
// NAND4 14
// AND8 1
// NAND3 1

module top (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
                  N430,N431,N432,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
        keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
                  keyinput125, keyinput126, keyinput127,
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
                  keyinput198, keyinput199,
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
        keyinput235);

  input keyinput200, keyinput201, keyinput202, keyinput203, keyinput204;
  input keyinput205, keyinput206, keyinput207, keyinput208, keyinput209;
  input keyinput210, keyinput211, keyinput212, keyinput213, keyinput214;
  input keyinput215, keyinput216, keyinput217, keyinput218, keyinput219;
  input keyinput220, keyinput221, keyinput222, keyinput223, keyinput224;
  input keyinput225, keyinput226, keyinput227, keyinput228, keyinput229;
  input keyinput230, keyinput231, keyinput232, keyinput233, keyinput234;
  input keyinput235;


  input keyinput128, keyinput129, keyinput130, keyinput131, keyinput132;
  input keyinput133, keyinput134, keyinput135, keyinput136, keyinput137;
  input keyinput138, keyinput139, keyinput140, keyinput141, keyinput142;
  input keyinput143, keyinput144, keyinput145, keyinput146, keyinput147;
  input keyinput148, keyinput149, keyinput150, keyinput151, keyinput152;
  input keyinput153, keyinput154, keyinput155, keyinput156, keyinput157;
  input keyinput158, keyinput159, keyinput160, keyinput161, keyinput162;
  input keyinput163, keyinput164, keyinput165, keyinput166, keyinput167;
  input keyinput168, keyinput169, keyinput170, keyinput171, keyinput172;
  input keyinput173, keyinput174, keyinput175, keyinput176, keyinput177;
  input keyinput178, keyinput179, keyinput180, keyinput181, keyinput182;
  input keyinput183, keyinput184, keyinput185, keyinput186, keyinput187;
  input keyinput188, keyinput189, keyinput190, keyinput191, keyinput192;
  input keyinput193, keyinput194, keyinput195, keyinput196, keyinput197;
  input keyinput198, keyinput199;

  wire KeyWire_0_1 , KeyWire_0_2;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31, keyinput32, keyinput33, keyinput34;
  input keyinput35, keyinput36, keyinput37, keyinput38, keyinput39;
  input keyinput40, keyinput41, keyinput42, keyinput43, keyinput44;
  input keyinput45, keyinput46, keyinput47, keyinput48, keyinput49;
  input keyinput50, keyinput51, keyinput52, keyinput53, keyinput54;
  input keyinput55, keyinput56, keyinput57, keyinput58, keyinput59;
  input keyinput60, keyinput61, keyinput62, keyinput63, keyinput64;
  input keyinput65, keyinput66, keyinput67, keyinput68, keyinput69;
  input keyinput70, keyinput71, keyinput72, keyinput73, keyinput74;
  input keyinput75, keyinput76, keyinput77, keyinput78, keyinput79;
  input keyinput80, keyinput81, keyinput82, keyinput83, keyinput84;
  input keyinput85, keyinput86, keyinput87, keyinput88, keyinput89;
  input keyinput90, keyinput91, keyinput92, keyinput93, keyinput94;
  input keyinput95, keyinput96, keyinput97, keyinput98, keyinput99;
  input keyinput100, keyinput101, keyinput102, keyinput103, keyinput104;
  input keyinput105, keyinput106, keyinput107, keyinput108, keyinput109;
  input keyinput110, keyinput111, keyinput112, keyinput113, keyinput114;
  input keyinput115, keyinput116, keyinput117, keyinput118, keyinput119;
  input keyinput120, keyinput121, keyinput122, keyinput123, keyinput124;
  input keyinput125, keyinput126, keyinput127;

  wire [0:127] keyinput_Wire_0;
  wire [0:64] KeyNOTWire_0;

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;

output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429;

  not NOT1_1 (keyinput_Wire_0[0], N1);
  xnor keyGate_0_0(N118, keyinput0, keyinput_Wire_0[0]);
  not NOT1_2 (keyinput_Wire_0[1], N4);
  xnor keyGate_0_1(KeyNOTWire_0[0], keyinput1, keyinput_Wire_0[1]);
  not KeyNOTGate_0_0(N119, KeyNOTWire_0[0]);
  not NOT1_3 (keyinput_Wire_0[2], N11);
  xnor keyGate_0_2(N122, keyinput2, keyinput_Wire_0[2]);
  not NOT1_4 (keyinput_Wire_0[3], N17);
  xnor keyGate_0_3(KeyNOTWire_0[1], keyinput3, keyinput_Wire_0[3]);
  not KeyNOTGate_0_1(N123, KeyNOTWire_0[1]);
  not NOT1_5 (keyinput_Wire_0[4], N24);
  xor keyGate_0_4(N126, keyinput4, keyinput_Wire_0[4]);
  not NOT1_6 (keyinput_Wire_0[5], N30);
  xor keyGate_0_5(KeyNOTWire_0[2], keyinput5, keyinput_Wire_0[5]);
  not KeyNOTGate_0_2(N127, KeyNOTWire_0[2]);
  not NOT1_7 (keyinput_Wire_0[6], N37);
  xnor keyGate_0_6(N130, keyinput6, keyinput_Wire_0[6]);
  not NOT1_8 (keyinput_Wire_0[7], N43);
  xor keyGate_0_7(N131, keyinput7, keyinput_Wire_0[7]);
  not NOT1_9 (keyinput_Wire_0[8], N50);
  xor keyGate_0_8(N134, keyinput8, keyinput_Wire_0[8]);
  not NOT1_10 (keyinput_Wire_0[9], N56);
  xnor keyGate_0_9(N135, keyinput9, keyinput_Wire_0[9]);
  not NOT1_11 (keyinput_Wire_0[10], N63);
  xnor keyGate_0_10(N138, keyinput10, keyinput_Wire_0[10]);
  not NOT1_12 (keyinput_Wire_0[11], N69);
  xor keyGate_0_11(KeyNOTWire_0[3], keyinput11, keyinput_Wire_0[11]);
  not KeyNOTGate_0_3(N139, KeyNOTWire_0[3]);
  not NOT1_13 (keyinput_Wire_0[12], N76);
  xnor keyGate_0_12(KeyNOTWire_0[4], keyinput12, keyinput_Wire_0[12]);
  not KeyNOTGate_0_4(N142, KeyNOTWire_0[4]);
  not NOT1_14 (keyinput_Wire_0[13], N82);
  xnor keyGate_0_13(N143, keyinput13, keyinput_Wire_0[13]);
  not NOT1_15 (keyinput_Wire_0[14], N89);
  xnor keyGate_0_14(N146, keyinput14, keyinput_Wire_0[14]);
  not NOT1_16 (keyinput_Wire_0[15], N95);
  xor keyGate_0_15(N147, keyinput15, keyinput_Wire_0[15]);
  not NOT1_17 (keyinput_Wire_0[16], N102);
  xor keyGate_0_16(KeyNOTWire_0[5], keyinput16, keyinput_Wire_0[16]);
  not KeyNOTGate_0_5(N150, KeyNOTWire_0[5]);
  not NOT1_18 (keyinput_Wire_0[17], N108);
  xor keyGate_0_17(N151, keyinput17, keyinput_Wire_0[17]);
  nand NAND2_19 (keyinput_Wire_0[18], N118, N4);
  xor keyGate_0_18(KeyNOTWire_0[6], keyinput18, keyinput_Wire_0[18]);
  not KeyNOTGate_0_6(N154, KeyNOTWire_0[6]);
  nor NOR2_20 (keyinput_Wire_0[19], N8, N119);
  xor keyGate_0_19(KeyNOTWire_0[7], keyinput19, keyinput_Wire_0[19]);
  not KeyNOTGate_0_7(N157, KeyNOTWire_0[7]);
nor NOR2_21 (N158, N14, N119);
  nand NAND2_22 (keyinput_Wire_0[20], N122, N17);
  xnor keyGate_0_20(N159, keyinput20, keyinput_Wire_0[20]);
  nand NAND2_23 (keyinput_Wire_0[21], N126, N30);
  xnor keyGate_0_21(KeyNOTWire_0[8], keyinput21, keyinput_Wire_0[21]);
  not KeyNOTGate_0_8(N162, KeyNOTWire_0[8]);
  nand NAND2_24 (keyinput_Wire_0[22], N130, N43);
  xor keyGate_0_22(KeyNOTWire_0[9], keyinput22, keyinput_Wire_0[22]);
  not KeyNOTGate_0_9(N165, KeyNOTWire_0[9]);
  nand NAND2_25 (keyinput_Wire_0[23], N134, N56);
  xnor keyGate_0_23(KeyNOTWire_0[10], keyinput23, keyinput_Wire_0[23]);
  not KeyNOTGate_0_10(N168, KeyNOTWire_0[10]);
  nand NAND2_26 (keyinput_Wire_0[24], N138, N69);
  xnor keyGate_0_24(N171, keyinput24, keyinput_Wire_0[24]);
  nand NAND2_27 (keyinput_Wire_0[25], N142, N82);
  xnor keyGate_0_25(KeyNOTWire_0[11], keyinput25, keyinput_Wire_0[25]);
  not KeyNOTGate_0_11(N174, KeyNOTWire_0[11]);
  nand NAND2_28 (keyinput_Wire_0[26], N146, N95);
  xor keyGate_0_26(KeyNOTWire_0[12], keyinput26, keyinput_Wire_0[26]);
  not KeyNOTGate_0_12(N177, KeyNOTWire_0[12]);
  nand NAND2_29 (keyinput_Wire_0[27], N150, N108);
  xor keyGate_0_27(N180, keyinput27, keyinput_Wire_0[27]);
  nor NOR2_30 (keyinput_Wire_0[28], N21, N123);
  xor keyGate_0_28(N183, keyinput28, keyinput_Wire_0[28]);
nor NOR2_31 (N184, N27, N123);
  nor NOR2_32 (keyinput_Wire_0[29], N34, N127);
  xnor keyGate_0_29(KeyNOTWire_0[13], keyinput29, keyinput_Wire_0[29]);
  not KeyNOTGate_0_13(N185, KeyNOTWire_0[13]);
nor NOR2_33 (N186, N40, N127);
  nor NOR2_34 (keyinput_Wire_0[30], N47, N131);
  xor keyGate_0_30(KeyNOTWire_0[14], keyinput30, keyinput_Wire_0[30]);
  not KeyNOTGate_0_14(N187, KeyNOTWire_0[14]);
nor NOR2_35 (N188, N53, N131);
  nor NOR2_36 (keyinput_Wire_0[31], N60, N135);
  xor keyGate_0_31(N189, keyinput31, keyinput_Wire_0[31]);
nor NOR2_37 (N190, N66, N135);
  nor NOR2_38 (keyinput_Wire_0[32], N73, N139);
  xnor keyGate_0_32(N191, keyinput32, keyinput_Wire_0[32]);
nor NOR2_39 (N192, N79, N139);
  nor NOR2_40 (keyinput_Wire_0[33], N86, N143);
  xor keyGate_0_33(KeyNOTWire_0[15], keyinput33, keyinput_Wire_0[33]);
  not KeyNOTGate_0_15(N193, KeyNOTWire_0[15]);
nor NOR2_41 (N194, N92, N143);
  nor NOR2_42 (keyinput_Wire_0[34], N99, N147);
  xnor keyGate_0_34(KeyNOTWire_0[16], keyinput34, keyinput_Wire_0[34]);
  not KeyNOTGate_0_16(N195, KeyNOTWire_0[16]);
nor NOR2_43 (N196, N105, N147);
  nor NOR2_44 (keyinput_Wire_0[35], N112, N151);
  xor keyGate_0_35(KeyNOTWire_0[17], keyinput35, keyinput_Wire_0[35]);
  not KeyNOTGate_0_17(N197, KeyNOTWire_0[17]);
nor NOR2_45 (N198, N115, N151);
  and AND9_46 (keyinput_Wire_0[36], N154, N159, N162, N165, N168, N171, N174, N177, N180);
  xnor keyGate_0_36(KeyNOTWire_0[18], keyinput36, keyinput_Wire_0[36]);
  not KeyNOTGate_0_18(N199, KeyNOTWire_0[18]);
  not NOT1_47 (keyinput_Wire_0[37], N199);
  xor keyGate_0_37(KeyNOTWire_0[19], keyinput37, keyinput_Wire_0[37]);
  not KeyNOTGate_0_19(N203, KeyNOTWire_0[19]);
not NOT1_48 (N213, N199);
not NOT1_49 (N223, N199);
  xor XOR2_50 (keyinput_Wire_0[38], N203, N154);
  xor keyGate_0_38(KeyNOTWire_0[20], keyinput38, keyinput_Wire_0[38]);
  not KeyNOTGate_0_20(N224, KeyNOTWire_0[20]);
  xor XOR2_51 (keyinput_Wire_0[39], N203, N159);
  xnor keyGate_0_39(N227, keyinput39, keyinput_Wire_0[39]);
  xor XOR2_52 (keyinput_Wire_0[40], N203, N162);
  xor keyGate_0_40(N230, keyinput40, keyinput_Wire_0[40]);
  xor XOR2_53 (keyinput_Wire_0[41], N203, N165);
  xor keyGate_0_41(N233, keyinput41, keyinput_Wire_0[41]);
  xor XOR2_54 (keyinput_Wire_0[42], N203, N168);
  xnor keyGate_0_42(N236, keyinput42, keyinput_Wire_0[42]);
  xor XOR2_55 (keyinput_Wire_0[43], N203, N171);
  xnor keyGate_0_43(N239, keyinput43, keyinput_Wire_0[43]);
nand NAND2_56 (N242, N1, N213);
  xor XOR2_57 (keyinput_Wire_0[44], N203, N174);
  xnor keyGate_0_44(KeyNOTWire_0[21], keyinput44, keyinput_Wire_0[44]);
  not KeyNOTGate_0_21(N243, KeyNOTWire_0[21]);
nand NAND2_58 (N246, N213, N11);
  xor XOR2_59 (keyinput_Wire_0[45], N203, N177);
  xnor keyGate_0_45(N247, keyinput45, keyinput_Wire_0[45]);
nand NAND2_60 (N250, N213, N24);
  xor XOR2_61 (keyinput_Wire_0[46], N203, N180);
  xor keyGate_0_46(KeyNOTWire_0[22], keyinput46, keyinput_Wire_0[46]);
  not KeyNOTGate_0_22(N251, KeyNOTWire_0[22]);
nand NAND2_62 (N254, N213, N37);
nand NAND2_63 (N255, N213, N50);
nand NAND2_64 (N256, N213, N63);
nand NAND2_65 (N257, N213, N76);
nand NAND2_66 (N258, N213, N89);
nand NAND2_67 (N259, N213, N102);
  nand NAND2_68 (keyinput_Wire_0[47], N224, N157);
  xnor keyGate_0_47(KeyNOTWire_0[23], keyinput47, keyinput_Wire_0[47]);
  not KeyNOTGate_0_23(N260, KeyNOTWire_0[23]);
  nand NAND2_69 (keyinput_Wire_0[48], N224, N158);
  xor keyGate_0_48(KeyNOTWire_0[24], keyinput48, keyinput_Wire_0[48]);
  not KeyNOTGate_0_24(N263, KeyNOTWire_0[24]);
  nand NAND2_70 (keyinput_Wire_0[49], N227, N183);
  xor keyGate_0_49(KeyNOTWire_0[25], keyinput49, keyinput_Wire_0[49]);
  not KeyNOTGate_0_25(N264, KeyNOTWire_0[25]);
  nand NAND2_71 (keyinput_Wire_0[50], N230, N185);
  xor keyGate_0_50(N267, keyinput50, keyinput_Wire_0[50]);
  nand NAND2_72 (keyinput_Wire_0[51], N233, N187);
  xnor keyGate_0_51(KeyNOTWire_0[26], keyinput51, keyinput_Wire_0[51]);
  not KeyNOTGate_0_26(N270, KeyNOTWire_0[26]);
  nand NAND2_73 (keyinput_Wire_0[52], N236, N189);
  xor keyGate_0_52(N273, keyinput52, keyinput_Wire_0[52]);
  nand NAND2_74 (keyinput_Wire_0[53], N239, N191);
  xnor keyGate_0_53(KeyNOTWire_0[27], keyinput53, keyinput_Wire_0[53]);
  not KeyNOTGate_0_27(N276, KeyNOTWire_0[27]);
  nand NAND2_75 (keyinput_Wire_0[54], N243, N193);
  xor keyGate_0_54(N279, keyinput54, keyinput_Wire_0[54]);
  nand NAND2_76 (keyinput_Wire_0[55], N247, N195);
  xor keyGate_0_55(KeyNOTWire_0[28], keyinput55, keyinput_Wire_0[55]);
  not KeyNOTGate_0_28(N282, KeyNOTWire_0[28]);
  nand NAND2_77 (keyinput_Wire_0[56], N251, N197);
  xor keyGate_0_56(KeyNOTWire_0[29], keyinput56, keyinput_Wire_0[56]);
  not KeyNOTGate_0_29(N285, KeyNOTWire_0[29]);
  nand NAND2_78 (keyinput_Wire_0[57], N227, N184);
  xnor keyGate_0_57(KeyNOTWire_0[30], keyinput57, keyinput_Wire_0[57]);
  not KeyNOTGate_0_30(N288, KeyNOTWire_0[30]);
  nand NAND2_79 (keyinput_Wire_0[58], N230, N186);
  xnor keyGate_0_58(KeyNOTWire_0[31], keyinput58, keyinput_Wire_0[58]);
  not KeyNOTGate_0_31(N289, KeyNOTWire_0[31]);
  nand NAND2_80 (keyinput_Wire_0[59], N233, N188);
  xnor keyGate_0_59(N290, keyinput59, keyinput_Wire_0[59]);
  nand NAND2_81 (keyinput_Wire_0[60], N236, N190);
  xor keyGate_0_60(KeyNOTWire_0[32], keyinput60, keyinput_Wire_0[60]);
  not KeyNOTGate_0_32(N291, KeyNOTWire_0[32]);
  nand NAND2_82 (keyinput_Wire_0[61], N239, N192);
  xnor keyGate_0_61(N292, keyinput61, keyinput_Wire_0[61]);
  nand NAND2_83 (keyinput_Wire_0[62], N243, N194);
  xnor keyGate_0_62(N293, keyinput62, keyinput_Wire_0[62]);
  nand NAND2_84 (keyinput_Wire_0[63], N247, N196);
  xnor keyGate_0_63(KeyNOTWire_0[33], keyinput63, keyinput_Wire_0[63]);
  not KeyNOTGate_0_33(N294, KeyNOTWire_0[33]);
  nand NAND2_85 (keyinput_Wire_0[64], N251, N198);
  xnor keyGate_0_64(N295, keyinput64, keyinput_Wire_0[64]);
  and AND9_86 (keyinput_Wire_0[65], N260, N264, N267, N270, N273, N276, N279, N282, N285);
  xor keyGate_0_65(KeyNOTWire_0[34], keyinput65, keyinput_Wire_0[65]);
  not KeyNOTGate_0_34(N296, KeyNOTWire_0[34]);
not NOT1_87 (N300, N263);
not NOT1_88 (N301, N288);
not NOT1_89 (N302, N289);
  not NOT1_90 (keyinput_Wire_0[66], N290);
  xor keyGate_0_66(N303, keyinput66, keyinput_Wire_0[66]);
  not NOT1_91 (keyinput_Wire_0[67], N291);
  xnor keyGate_0_67(KeyNOTWire_0[35], keyinput67, keyinput_Wire_0[67]);
  not KeyNOTGate_0_35(N304, KeyNOTWire_0[35]);
  not NOT1_92 (keyinput_Wire_0[68], N292);
  xor keyGate_0_68(KeyNOTWire_0[36], keyinput68, keyinput_Wire_0[68]);
  not KeyNOTGate_0_36(N305, KeyNOTWire_0[36]);
  not NOT1_93 (keyinput_Wire_0[69], N293);
  xnor keyGate_0_69(N306, keyinput69, keyinput_Wire_0[69]);
not NOT1_94 (N307, N294);
  not NOT1_95 (keyinput_Wire_0[70], N295);
  xnor keyGate_0_70(KeyNOTWire_0[37], keyinput70, keyinput_Wire_0[70]);
  not KeyNOTGate_0_37(N308, KeyNOTWire_0[37]);
  not NOT1_96 (keyinput_Wire_0[71], N296);
  xor keyGate_0_71(N309, keyinput71, keyinput_Wire_0[71]);
  not NOT1_97 (keyinput_Wire_0[72], N296);
  xnor keyGate_0_72(N319, keyinput72, keyinput_Wire_0[72]);
not NOT1_98 (KeyWire_0_1, N296);
  xor flip_it (N329, KeyWire_0_1, KeyWire_0_2 );
  xor XOR2_99 (keyinput_Wire_0[73], N309, N260);
  xor keyGate_0_73(N330, keyinput73, keyinput_Wire_0[73]);
  xor XOR2_100 (keyinput_Wire_0[74], N309, N264);
  xor keyGate_0_74(N331, keyinput74, keyinput_Wire_0[74]);
  xor XOR2_101 (keyinput_Wire_0[75], N309, N267);
  xnor keyGate_0_75(KeyNOTWire_0[38], keyinput75, keyinput_Wire_0[75]);
  not KeyNOTGate_0_38(N332, KeyNOTWire_0[38]);
  xor XOR2_102 (keyinput_Wire_0[76], N309, N270);
  xnor keyGate_0_76(N333, keyinput76, keyinput_Wire_0[76]);
nand NAND2_103 (N334, N8, N319);
  xor XOR2_104 (keyinput_Wire_0[77], N309, N273);
  xnor keyGate_0_77(N335, keyinput77, keyinput_Wire_0[77]);
nand NAND2_105 (N336, N319, N21);
  xor XOR2_106 (keyinput_Wire_0[78], N309, N276);
  xnor keyGate_0_78(KeyNOTWire_0[39], keyinput78, keyinput_Wire_0[78]);
  not KeyNOTGate_0_39(N337, KeyNOTWire_0[39]);
  nand NAND2_107 (keyinput_Wire_0[79], N319, N34);
  xnor keyGate_0_79(KeyNOTWire_0[40], keyinput79, keyinput_Wire_0[79]);
  not KeyNOTGate_0_40(N338, KeyNOTWire_0[40]);
  xor XOR2_108 (keyinput_Wire_0[80], N309, N279);
  xor keyGate_0_80(KeyNOTWire_0[41], keyinput80, keyinput_Wire_0[80]);
  not KeyNOTGate_0_41(N339, KeyNOTWire_0[41]);
  nand NAND2_109 (keyinput_Wire_0[81], N319, N47);
  xnor keyGate_0_81(N340, keyinput81, keyinput_Wire_0[81]);
  xor XOR2_110 (keyinput_Wire_0[82], N309, N282);
  xnor keyGate_0_82(N341, keyinput82, keyinput_Wire_0[82]);
nand NAND2_111 (N342, N319, N60);
  xor XOR2_112 (keyinput_Wire_0[83], N309, N285);
  xor keyGate_0_83(N343, keyinput83, keyinput_Wire_0[83]);
nand NAND2_113 (N344, N319, N73);
nand NAND2_114 (N345, N319, N86);
nand NAND2_115 (N346, N319, N99);
nand NAND2_116 (N347, N319, N112);
  nand NAND2_117 (keyinput_Wire_0[84], N330, N300);
  xor keyGate_0_84(N348, keyinput84, keyinput_Wire_0[84]);
  nand NAND2_118 (keyinput_Wire_0[85], N331, N301);
  xnor keyGate_0_85(N349, keyinput85, keyinput_Wire_0[85]);
  nand NAND2_119 (keyinput_Wire_0[86], N332, N302);
  xor keyGate_0_86(KeyNOTWire_0[42], keyinput86, keyinput_Wire_0[86]);
  not KeyNOTGate_0_42(N350, KeyNOTWire_0[42]);
  nand NAND2_120 (keyinput_Wire_0[87], N333, N303);
  xnor keyGate_0_87(N351, keyinput87, keyinput_Wire_0[87]);
  nand NAND2_121 (keyinput_Wire_0[88], N335, N304);
  xnor keyGate_0_88(KeyNOTWire_0[43], keyinput88, keyinput_Wire_0[88]);
  not KeyNOTGate_0_43(N352, KeyNOTWire_0[43]);
  nand NAND2_122 (keyinput_Wire_0[89], N337, N305);
  xor keyGate_0_89(N353, keyinput89, keyinput_Wire_0[89]);
  nand NAND2_123 (keyinput_Wire_0[90], N339, N306);
  xnor keyGate_0_90(KeyNOTWire_0[44], keyinput90, keyinput_Wire_0[90]);
  not KeyNOTGate_0_44(N354, KeyNOTWire_0[44]);
  nand NAND2_124 (keyinput_Wire_0[91], N341, N307);
  xnor keyGate_0_91(N355, keyinput91, keyinput_Wire_0[91]);
  nand NAND2_125 (keyinput_Wire_0[92], N343, N308);
  xnor keyGate_0_92(KeyNOTWire_0[45], keyinput92, keyinput_Wire_0[92]);
  not KeyNOTGate_0_45(N356, KeyNOTWire_0[45]);
  and AND9_126 (keyinput_Wire_0[93], N348, N349, N350, N351, N352, N353, N354, N355, N356);
  xor keyGate_0_93(N357, keyinput93, keyinput_Wire_0[93]);
  not NOT1_127 (keyinput_Wire_0[94], N357);
  xor keyGate_0_94(N360, keyinput94, keyinput_Wire_0[94]);
  not NOT1_128 (keyinput_Wire_0[95], N357);
  xor keyGate_0_95(KeyNOTWire_0[46], keyinput95, keyinput_Wire_0[95]);
  not KeyNOTGate_0_46(N370, KeyNOTWire_0[46]);
  nand NAND2_129 (keyinput_Wire_0[96], N14, N360);
  xnor keyGate_0_96(N371, keyinput96, keyinput_Wire_0[96]);
  nand NAND2_130 (keyinput_Wire_0[97], N360, N27);
  xor keyGate_0_97(KeyNOTWire_0[47], keyinput97, keyinput_Wire_0[97]);
  not KeyNOTGate_0_47(N372, KeyNOTWire_0[47]);
  nand NAND2_131 (keyinput_Wire_0[98], N360, N40);
  xor keyGate_0_98(KeyNOTWire_0[48], keyinput98, keyinput_Wire_0[98]);
  not KeyNOTGate_0_48(N373, KeyNOTWire_0[48]);
  nand NAND2_132 (keyinput_Wire_0[99], N360, N53);
  xor keyGate_0_99(KeyNOTWire_0[49], keyinput99, keyinput_Wire_0[99]);
  not KeyNOTGate_0_49(N374, KeyNOTWire_0[49]);
  nand NAND2_133 (keyinput_Wire_0[100], N360, N66);
  xor keyGate_0_100(KeyNOTWire_0[50], keyinput100, keyinput_Wire_0[100]);
  not KeyNOTGate_0_50(N375, KeyNOTWire_0[50]);
  nand NAND2_134 (keyinput_Wire_0[101], N360, N79);
  xor keyGate_0_101(N376, keyinput101, keyinput_Wire_0[101]);
  nand NAND2_135 (keyinput_Wire_0[102], N360, N92);
  xor keyGate_0_102(KeyNOTWire_0[51], keyinput102, keyinput_Wire_0[102]);
  not KeyNOTGate_0_51(N377, KeyNOTWire_0[51]);
  nand NAND2_136 (keyinput_Wire_0[103], N360, N105);
  xor keyGate_0_103(KeyNOTWire_0[52], keyinput103, keyinput_Wire_0[103]);
  not KeyNOTGate_0_52(N378, KeyNOTWire_0[52]);
  nand NAND2_137 (keyinput_Wire_0[104], N360, N115);
  xnor keyGate_0_104(KeyNOTWire_0[53], keyinput104, keyinput_Wire_0[104]);
  not KeyNOTGate_0_53(N379, KeyNOTWire_0[53]);
  nand NAND4_138 (keyinput_Wire_0[105], N4, N242, N334, N371);
  xor keyGate_0_105(N380, keyinput105, keyinput_Wire_0[105]);
  nand NAND4_139 (keyinput_Wire_0[106], N246, N336, N372, N17);
  xnor keyGate_0_106(N381, keyinput106, keyinput_Wire_0[106]);
  nand NAND4_140 (keyinput_Wire_0[107], N250, N338, N373, N30);
  xnor keyGate_0_107(KeyNOTWire_0[54], keyinput107, keyinput_Wire_0[107]);
  not KeyNOTGate_0_54(N386, KeyNOTWire_0[54]);
  nand NAND4_141 (keyinput_Wire_0[108], N254, N340, N374, N43);
  xnor keyGate_0_108(KeyNOTWire_0[55], keyinput108, keyinput_Wire_0[108]);
  not KeyNOTGate_0_55(N393, KeyNOTWire_0[55]);
  nand NAND4_142 (keyinput_Wire_0[109], N255, N342, N375, N56);
  xor keyGate_0_109(N399, keyinput109, keyinput_Wire_0[109]);
  nand NAND4_143 (keyinput_Wire_0[110], N256, N344, N376, N69);
  xnor keyGate_0_110(KeyNOTWire_0[56], keyinput110, keyinput_Wire_0[110]);
  not KeyNOTGate_0_56(N404, KeyNOTWire_0[56]);
  nand NAND4_144 (keyinput_Wire_0[111], N257, N345, N377, N82);
  xnor keyGate_0_111(KeyNOTWire_0[57], keyinput111, keyinput_Wire_0[111]);
  not KeyNOTGate_0_57(N407, KeyNOTWire_0[57]);
  nand NAND4_145 (keyinput_Wire_0[112], N258, N346, N378, N95);
  xor keyGate_0_112(KeyNOTWire_0[58], keyinput112, keyinput_Wire_0[112]);
  not KeyNOTGate_0_58(N411, KeyNOTWire_0[58]);
  nand NAND4_146 (keyinput_Wire_0[113], N259, N347, N379, N108);
  xor keyGate_0_113(N414, keyinput113, keyinput_Wire_0[113]);
  not NOT1_147 (keyinput_Wire_0[114], N380);
  xor keyGate_0_114(N415, keyinput114, keyinput_Wire_0[114]);
  and AND8_148 (keyinput_Wire_0[115], N381, N386, N393, N399, N404, N407, N411, N414);
  xnor keyGate_0_115(KeyNOTWire_0[59], keyinput115, keyinput_Wire_0[115]);
  not KeyNOTGate_0_59(N416, KeyNOTWire_0[59]);
  not NOT1_149 (keyinput_Wire_0[116], N393);
  xnor keyGate_0_116(N417, keyinput116, keyinput_Wire_0[116]);
  not NOT1_150 (keyinput_Wire_0[117], N404);
  xor keyGate_0_117(KeyNOTWire_0[60], keyinput117, keyinput_Wire_0[117]);
  not KeyNOTGate_0_60(N418, KeyNOTWire_0[60]);
  not NOT1_151 (keyinput_Wire_0[118], N407);
  xnor keyGate_0_118(KeyNOTWire_0[61], keyinput118, keyinput_Wire_0[118]);
  not KeyNOTGate_0_61(N419, KeyNOTWire_0[61]);
  not NOT1_152 (keyinput_Wire_0[119], N411);
  xor keyGate_0_119(N420, keyinput119, keyinput_Wire_0[119]);
  nor NOR2_153 (keyinput_Wire_0[120], N415, N416);
  xor keyGate_0_120(KeyNOTWire_0[62], keyinput120, keyinput_Wire_0[120]);
  not KeyNOTGate_0_62(N421, KeyNOTWire_0[62]);
  nand NAND2_154 (keyinput_Wire_0[121], N386, N417);
  xnor keyGate_0_121(KeyNOTWire_0[63], keyinput121, keyinput_Wire_0[121]);
  not KeyNOTGate_0_63(N422, KeyNOTWire_0[63]);
  nand NAND4_155 (keyinput_Wire_0[122], N386, N393, N418, N399);
  xor keyGate_0_122(N425, keyinput122, keyinput_Wire_0[122]);
  nand NAND3_156 (keyinput_Wire_0[123], N399, N393, N419);
  xnor keyGate_0_123(N428, keyinput123, keyinput_Wire_0[123]);
  nand NAND4_157 (keyinput_Wire_0[124], N386, N393, N407, N420);
  xnor keyGate_0_124(N429, keyinput124, keyinput_Wire_0[124]);
  nand NAND4_158 (keyinput_Wire_0[125], N381, N386, N422, N399);
  xnor keyGate_0_125(N430, keyinput125, keyinput_Wire_0[125]);
  nand NAND4_159 (keyinput_Wire_0[126], N381, N386, N425, N428);
  xnor keyGate_0_126(N431, keyinput126, keyinput_Wire_0[126]);
  nand NAND4_160 (keyinput_Wire_0[127], N381, N422, N425, N429);
  xor keyGate_0_127(KeyNOTWire_0[64], keyinput127, keyinput_Wire_0[127]);
  not KeyNOTGate_0_64(N432, KeyNOTWire_0[64]);

AntiSAT some_name( KeyWire_0_2, N8, N4, N99, N76, N21, N66, N17, N73, N34, N50, N43, N47, N95, N79, N108, N1, N60, N92, N56, N40, N105, N102, N86, N115, N112, N30, N24, N69, N89, N53, N37, N11, N82, N63, N14, N27, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
       keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
       keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
       keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
       keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
       keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
       keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
       keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
       keyinput235);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N8, N4, N99, N76, N21, N66, N17, N73, N34, N50, N43, N47, N95, N79, N108, N1, N60, N92, N56, N40, N105, N102, N86, N115, N112, N30, N24, N69, N89, N53, N37, N11, N82, N63, N14, N27, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199 ,
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
        keyinput235);

  input keyinput200, keyinput201, keyinput202, keyinput203, keyinput204;
  input keyinput205, keyinput206, keyinput207, keyinput208, keyinput209;
  input keyinput210, keyinput211, keyinput212, keyinput213, keyinput214;
  input keyinput215, keyinput216, keyinput217, keyinput218, keyinput219;
  input keyinput220, keyinput221, keyinput222, keyinput223, keyinput224;
  input keyinput225, keyinput226, keyinput227, keyinput228, keyinput229;
  input keyinput230, keyinput231, keyinput232, keyinput233, keyinput234;
  input keyinput235;

  wire [0:35] keyNTin_Wire_1;
  wire [0:13] KeyNOTWire_1;

  input N8, N4, N99, N76, N21, N66, N17, N73, N34, N50, N43, N47, N95, N79, N108, N1, N60, N92, N56, N40, N105, N102, N86, N115, N112, N30, N24, N69, N89, N53, N37, N11, N82, N63, N14, N27;
  input keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73 ;

  xnor KeyGate0 (newWire_0, N8, keyinput128);
  xnor KeyGate1 (newWire_1, N4, keyinput129);
  xnor KeyGate2 (newWire_2, N99, keyinput130);
  xor  KeyGate3 (keyNTin_Wire_1[0], N76, keyinput131);
  xnor keyNTinGate_1_0(newWire_3, keyinput200, keyNTin_Wire_1[0]);
  xor  KeyGate4 (newWire_4, N21, keyinput132);
  xnor KeyGate5 (keyNTin_Wire_1[1], N66, keyinput133);
  xnor keyNTinGate_1_1(newWire_5, keyinput201, keyNTin_Wire_1[1]);
  xor  KeyGate6 (newWire_6, N17, keyinput134);
  xor  KeyGate7 (keyNTin_Wire_1[2], N73, keyinput135);
  xor keyNTinGate_1_2(KeyNOTWire_1[0], keyinput202, keyNTin_Wire_1[2]);
  not KeyNOTGate_1_0(newWire_7, KeyNOTWire_1[0]);
  xnor KeyGate8 (keyNTin_Wire_1[3], N34, keyinput136);
  xor keyNTinGate_1_3(newWire_8, keyinput203, keyNTin_Wire_1[3]);
  xor  KeyGate9 (keyNTin_Wire_1[4], N50, keyinput137);
  xnor keyNTinGate_1_4(KeyNOTWire_1[1], keyinput204, keyNTin_Wire_1[4]);
  not KeyNOTGate_1_1(newWire_9, KeyNOTWire_1[1]);
  xor  KeyGate10 (keyNTin_Wire_1[5], N43, keyinput138);
  xor keyNTinGate_1_5(KeyNOTWire_1[2], keyinput205, keyNTin_Wire_1[5]);
  not KeyNOTGate_1_2(newWire_10, KeyNOTWire_1[2]);
  xor  KeyGate11 (keyNTin_Wire_1[6], N47, keyinput139);
  xnor keyNTinGate_1_6(KeyNOTWire_1[3], keyinput206, keyNTin_Wire_1[6]);
  not KeyNOTGate_1_3(newWire_11, KeyNOTWire_1[3]);
  xor  KeyGate12 (keyNTin_Wire_1[7], N95, keyinput140);
  xnor keyNTinGate_1_7(newWire_12, keyinput207, keyNTin_Wire_1[7]);
  xor  KeyGate13 (keyNTin_Wire_1[8], N79, keyinput141);
  xor keyNTinGate_1_8(newWire_13, keyinput208, keyNTin_Wire_1[8]);
  xnor KeyGate14 (keyNTin_Wire_1[9], N108, keyinput142);
  xnor keyNTinGate_1_9(newWire_14, keyinput209, keyNTin_Wire_1[9]);
  xnor KeyGate15 (keyNTin_Wire_1[10], N1, keyinput143);
  xnor keyNTinGate_1_10(newWire_15, keyinput210, keyNTin_Wire_1[10]);
  xor  KeyGate16 (keyNTin_Wire_1[11], N60, keyinput144);
  xnor keyNTinGate_1_11(KeyNOTWire_1[4], keyinput211, keyNTin_Wire_1[11]);
  not KeyNOTGate_1_4(newWire_16, KeyNOTWire_1[4]);
  xor  KeyGate17 (keyNTin_Wire_1[12], N92, keyinput145);
  xor keyNTinGate_1_12(newWire_17, keyinput212, keyNTin_Wire_1[12]);
  xor  KeyGate18 (newWire_18, N56, keyinput146);
  xor  KeyGate19 (keyNTin_Wire_1[13], N40, keyinput147);
  xor keyNTinGate_1_13(KeyNOTWire_1[5], keyinput213, keyNTin_Wire_1[13]);
  not KeyNOTGate_1_5(newWire_19, KeyNOTWire_1[5]);
  xor  KeyGate20 (newWire_20, N105, keyinput148);
  xnor KeyGate21 (newWire_21, N102, keyinput149);
  xnor KeyGate22 (keyNTin_Wire_1[14], N86, keyinput150);
  xor keyNTinGate_1_14(newWire_22, keyinput214, keyNTin_Wire_1[14]);
  xnor KeyGate23 (keyNTin_Wire_1[15], N115, keyinput151);
  xnor keyNTinGate_1_15(newWire_23, keyinput215, keyNTin_Wire_1[15]);
  xnor KeyGate24 (newWire_24, N112, keyinput152);
  xor  KeyGate25 (keyNTin_Wire_1[16], N30, keyinput153);
  xor keyNTinGate_1_16(newWire_25, keyinput216, keyNTin_Wire_1[16]);
  xor  KeyGate26 (keyNTin_Wire_1[17], N24, keyinput154);
  xnor keyNTinGate_1_17(newWire_26, keyinput217, keyNTin_Wire_1[17]);
  xor  KeyGate27 (newWire_27, N69, keyinput155);
  xor  KeyGate28 (newWire_28, N89, keyinput156);
  xor  KeyGate29 (newWire_29, N53, keyinput157);
  xnor KeyGate30 (newWire_30, N37, keyinput158);
  xnor KeyGate31 (newWire_31, N11, keyinput159);
  xnor KeyGate32 (newWire_32, N82, keyinput160);
  xnor KeyGate33 (keyNTin_Wire_1[18], N63, keyinput161);
  xor keyNTinGate_1_18(newWire_33, keyinput218, keyNTin_Wire_1[18]);
  xor  KeyGate34 (newWire_34, N14, keyinput162);
  xnor KeyGate35 (keyNTin_Wire_1[19], N27, keyinput163);
  xnor keyNTinGate_1_19(newWire_35, keyinput219, keyNTin_Wire_1[19]);
  xnor KeyGate36 (newWire_36, N8, keyinput164);
  xor  KeyGate37 (keyNTin_Wire_1[20], N4, keyinput165);
  xnor keyNTinGate_1_20(newWire_37, keyinput220, keyNTin_Wire_1[20]);
  xnor KeyGate38 (keyNTin_Wire_1[21], N99, keyinput166);
  xor keyNTinGate_1_21(newWire_38, keyinput221, keyNTin_Wire_1[21]);
  xnor KeyGate39 (newWire_39, N76, keyinput167);
  xnor KeyGate40 (keyNTin_Wire_1[22], N21, keyinput168);
  xor keyNTinGate_1_22(KeyNOTWire_1[6], keyinput222, keyNTin_Wire_1[22]);
  not KeyNOTGate_1_6(newWire_40, KeyNOTWire_1[6]);
  xnor KeyGate41 (newWire_41, N66, keyinput169);
  xnor KeyGate42 (keyNTin_Wire_1[23], N17, keyinput170);
  xor keyNTinGate_1_23(KeyNOTWire_1[7], keyinput223, keyNTin_Wire_1[23]);
  not KeyNOTGate_1_7(newWire_42, KeyNOTWire_1[7]);
  xnor KeyGate43 (newWire_43, N73, keyinput171);
  xnor KeyGate44 (newWire_44, N34, keyinput172);
  xor  KeyGate45 (keyNTin_Wire_1[24], N50, keyinput173);
  xor keyNTinGate_1_24(KeyNOTWire_1[8], keyinput224, keyNTin_Wire_1[24]);
  not KeyNOTGate_1_8(newWire_45, KeyNOTWire_1[8]);
  xnor KeyGate46 (newWire_46, N43, keyinput174);
  xor  KeyGate47 (keyNTin_Wire_1[25], N47, keyinput175);
  xor keyNTinGate_1_25(KeyNOTWire_1[9], keyinput225, keyNTin_Wire_1[25]);
  not KeyNOTGate_1_9(newWire_47, KeyNOTWire_1[9]);
  xnor KeyGate48 (keyNTin_Wire_1[26], N95, keyinput176);
  xor keyNTinGate_1_26(KeyNOTWire_1[10], keyinput226, keyNTin_Wire_1[26]);
  not KeyNOTGate_1_10(newWire_48, KeyNOTWire_1[10]);
  xor  KeyGate49 (newWire_49, N79, keyinput177);
  xor  KeyGate50 (newWire_50, N108, keyinput178);
  xor  KeyGate51 (keyNTin_Wire_1[27], N1, keyinput179);
  xnor keyNTinGate_1_27(newWire_51, keyinput227, keyNTin_Wire_1[27]);
  xor  KeyGate52 (newWire_52, N60, keyinput180);
  xor  KeyGate53 (newWire_53, N92, keyinput181);
  xor  KeyGate54 (keyNTin_Wire_1[28], N56, keyinput182);
  xnor keyNTinGate_1_28(newWire_54, keyinput228, keyNTin_Wire_1[28]);
  xnor KeyGate55 (newWire_55, N40, keyinput183);
  xor  KeyGate56 (newWire_56, N105, keyinput184);
  xor  KeyGate57 (newWire_57, N102, keyinput185);
  xor  KeyGate58 (newWire_58, N86, keyinput186);
  xnor KeyGate59 (newWire_59, N115, keyinput187);
  xnor KeyGate60 (newWire_60, N112, keyinput188);
  xor  KeyGate61 (keyNTin_Wire_1[29], N30, keyinput189);
  xor keyNTinGate_1_29(newWire_61, keyinput229, keyNTin_Wire_1[29]);
  xnor KeyGate62 (keyNTin_Wire_1[30], N24, keyinput190);
  xor keyNTinGate_1_30(KeyNOTWire_1[11], keyinput230, keyNTin_Wire_1[30]);
  not KeyNOTGate_1_11(newWire_62, KeyNOTWire_1[11]);
  xnor KeyGate63 (newWire_63, N69, keyinput191);
  xnor KeyGate64 (keyNTin_Wire_1[31], N89, keyinput192);
  xor keyNTinGate_1_31(KeyNOTWire_1[12], keyinput231, keyNTin_Wire_1[31]);
  not KeyNOTGate_1_12(newWire_64, KeyNOTWire_1[12]);
  xnor KeyGate65 (newWire_65, N53, keyinput193);
  xor  KeyGate66 (keyNTin_Wire_1[32], N37, keyinput194);
  xor keyNTinGate_1_32(newWire_66, keyinput232, keyNTin_Wire_1[32]);
  xnor KeyGate67 (keyNTin_Wire_1[33], N11, keyinput195);
  xnor keyNTinGate_1_33(newWire_67, keyinput233, keyNTin_Wire_1[33]);
  xor  KeyGate68 (keyNTin_Wire_1[34], N82, keyinput196);
  xor keyNTinGate_1_34(newWire_68, keyinput234, keyNTin_Wire_1[34]);
  xnor KeyGate69 (keyNTin_Wire_1[35], N63, keyinput197);
  xnor keyNTinGate_1_35(KeyNOTWire_1[13], keyinput235, keyNTin_Wire_1[35]);
  not KeyNOTGate_1_13(newWire_69, KeyNOTWire_1[13]);
  xor  KeyGate70 (newWire_70, N14, keyinput198);
  xnor KeyGate71 (newWire_71, N27, keyinput199);
  and some_function (newWire_72, newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35 );
  nand compl_function (newWire_73, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71);
  and finalAND (KeyWire_0_2, newWire_72, newWire_73);

endmodule /* AntiSAT */
