`timescale 1ns / 1ps
// Verilog
// c880
// Ninputs 60
// Noutputs 26
// NtotalGates 383
// NAND4 13
// AND3 12
// NAND2 60
// NAND3 14
// AND2 105
// OR2 29
// NOT1 63
// NOR2 61
// BUFF1 26

module top (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
                  N865,N866,N874,N878,N879,N880,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
        keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
        keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
        keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
        keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
        keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
        keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
        keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
        keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
        keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
        keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
        keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
        keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
        keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
        keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
        keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
        keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
        keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
                  keyinput255,
        keyinput256, keyinput257, keyinput258, keyinput259, keyinput260,
        keyinput261, keyinput262, keyinput263, keyinput264, keyinput265,
        keyinput266, keyinput267, keyinput268, keyinput269, keyinput270,
        keyinput271, keyinput272, keyinput273, keyinput274, keyinput275,
        keyinput276, keyinput277, keyinput278, keyinput279, keyinput280,
        keyinput281, keyinput282, keyinput283, keyinput284, keyinput285,
        keyinput286, keyinput287, keyinput288, keyinput289, keyinput290,
        keyinput291, keyinput292, keyinput293, keyinput294, keyinput295,
        keyinput296, keyinput297, keyinput298, keyinput299, keyinput300,
        keyinput301, keyinput302, keyinput303, keyinput304, keyinput305,
        keyinput306, keyinput307, keyinput308, keyinput309, keyinput310,
        keyinput311, keyinput312, keyinput313, keyinput314, keyinput315,
        keyinput316, keyinput317, keyinput318, keyinput319, keyinput320,
        keyinput321, keyinput322, keyinput323, keyinput324, keyinput325,
        keyinput326, keyinput327, keyinput328, keyinput329, keyinput330,
        keyinput331, keyinput332, keyinput333, keyinput334, keyinput335,
        keyinput336, keyinput337, keyinput338, keyinput339, keyinput340,
        keyinput341, keyinput342, keyinput343, keyinput344, keyinput345,
        keyinput346, keyinput347, keyinput348, keyinput349, keyinput350,
        keyinput351, keyinput352, keyinput353, keyinput354, keyinput355,
        keyinput356, keyinput357, keyinput358, keyinput359, keyinput360,
        keyinput361, keyinput362, keyinput363, keyinput364, keyinput365,
        keyinput366, keyinput367, keyinput368, keyinput369, keyinput370,
                  keyinput371, keyinput372, keyinput373, keyinput374, keyinput375,
        keyinput376, keyinput377, keyinput378, keyinput379, keyinput380,
        keyinput381, keyinput382, keyinput383, keyinput384, keyinput385,
        keyinput386, keyinput387, keyinput388, keyinput389, keyinput390,
        keyinput391, keyinput392, keyinput393, keyinput394, keyinput395,
        keyinput396, keyinput397, keyinput398, keyinput399, keyinput400,
        keyinput401, keyinput402, keyinput403, keyinput404, keyinput405,
        keyinput406, keyinput407, keyinput408, keyinput409, keyinput410,
        keyinput411, keyinput412, keyinput413, keyinput414, keyinput415,
        keyinput416, keyinput417, keyinput418, keyinput419, keyinput420,
        keyinput421, keyinput422, keyinput423, keyinput424, keyinput425,
        keyinput426, keyinput427, keyinput428, keyinput429, keyinput430,
        keyinput431, keyinput432, keyinput433, keyinput434, keyinput435);

  input keyinput376, keyinput377, keyinput378, keyinput379, keyinput380;
  input keyinput381, keyinput382, keyinput383, keyinput384, keyinput385;
  input keyinput386, keyinput387, keyinput388, keyinput389, keyinput390;
  input keyinput391, keyinput392, keyinput393, keyinput394, keyinput395;
  input keyinput396, keyinput397, keyinput398, keyinput399, keyinput400;
  input keyinput401, keyinput402, keyinput403, keyinput404, keyinput405;
  input keyinput406, keyinput407, keyinput408, keyinput409, keyinput410;
  input keyinput411, keyinput412, keyinput413, keyinput414, keyinput415;
  input keyinput416, keyinput417, keyinput418, keyinput419, keyinput420;
  input keyinput421, keyinput422, keyinput423, keyinput424, keyinput425;
  input keyinput426, keyinput427, keyinput428, keyinput429, keyinput430;
  input keyinput431, keyinput432, keyinput433, keyinput434, keyinput435;


  input keyinput256, keyinput257, keyinput258, keyinput259, keyinput260;
  input keyinput261, keyinput262, keyinput263, keyinput264, keyinput265;
  input keyinput266, keyinput267, keyinput268, keyinput269, keyinput270;
  input keyinput271, keyinput272, keyinput273, keyinput274, keyinput275;
  input keyinput276, keyinput277, keyinput278, keyinput279, keyinput280;
  input keyinput281, keyinput282, keyinput283, keyinput284, keyinput285;
  input keyinput286, keyinput287, keyinput288, keyinput289, keyinput290;
  input keyinput291, keyinput292, keyinput293, keyinput294, keyinput295;
  input keyinput296, keyinput297, keyinput298, keyinput299, keyinput300;
  input keyinput301, keyinput302, keyinput303, keyinput304, keyinput305;
  input keyinput306, keyinput307, keyinput308, keyinput309, keyinput310;
  input keyinput311, keyinput312, keyinput313, keyinput314, keyinput315;
  input keyinput316, keyinput317, keyinput318, keyinput319, keyinput320;
  input keyinput321, keyinput322, keyinput323, keyinput324, keyinput325;
  input keyinput326, keyinput327, keyinput328, keyinput329, keyinput330;
  input keyinput331, keyinput332, keyinput333, keyinput334, keyinput335;
  input keyinput336, keyinput337, keyinput338, keyinput339, keyinput340;
  input keyinput341, keyinput342, keyinput343, keyinput344, keyinput345;
  input keyinput346, keyinput347, keyinput348, keyinput349, keyinput350;
  input keyinput351, keyinput352, keyinput353, keyinput354, keyinput355;
  input keyinput356, keyinput357, keyinput358, keyinput359, keyinput360;
  input keyinput361, keyinput362, keyinput363, keyinput364, keyinput365;
  input keyinput366, keyinput367, keyinput368, keyinput369, keyinput370;
  input keyinput371, keyinput372, keyinput373, keyinput374, keyinput375;

  wire KeyWire_0_1 , KeyWire_0_2, keyinput_Wire_1;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31, keyinput32, keyinput33, keyinput34;
  input keyinput35, keyinput36, keyinput37, keyinput38, keyinput39;
  input keyinput40, keyinput41, keyinput42, keyinput43, keyinput44;
  input keyinput45, keyinput46, keyinput47, keyinput48, keyinput49;
  input keyinput50, keyinput51, keyinput52, keyinput53, keyinput54;
  input keyinput55, keyinput56, keyinput57, keyinput58, keyinput59;
  input keyinput60, keyinput61, keyinput62, keyinput63, keyinput64;
  input keyinput65, keyinput66, keyinput67, keyinput68, keyinput69;
  input keyinput70, keyinput71, keyinput72, keyinput73, keyinput74;
  input keyinput75, keyinput76, keyinput77, keyinput78, keyinput79;
  input keyinput80, keyinput81, keyinput82, keyinput83, keyinput84;
  input keyinput85, keyinput86, keyinput87, keyinput88, keyinput89;
  input keyinput90, keyinput91, keyinput92, keyinput93, keyinput94;
  input keyinput95, keyinput96, keyinput97, keyinput98, keyinput99;
  input keyinput100, keyinput101, keyinput102, keyinput103, keyinput104;
  input keyinput105, keyinput106, keyinput107, keyinput108, keyinput109;
  input keyinput110, keyinput111, keyinput112, keyinput113, keyinput114;
  input keyinput115, keyinput116, keyinput117, keyinput118, keyinput119;
  input keyinput120, keyinput121, keyinput122, keyinput123, keyinput124;
  input keyinput125, keyinput126, keyinput127, keyinput128, keyinput129;
  input keyinput130, keyinput131, keyinput132, keyinput133, keyinput134;
  input keyinput135, keyinput136, keyinput137, keyinput138, keyinput139;
  input keyinput140, keyinput141, keyinput142, keyinput143, keyinput144;
  input keyinput145, keyinput146, keyinput147, keyinput148, keyinput149;
  input keyinput150, keyinput151, keyinput152, keyinput153, keyinput154;
  input keyinput155, keyinput156, keyinput157, keyinput158, keyinput159;
  input keyinput160, keyinput161, keyinput162, keyinput163, keyinput164;
  input keyinput165, keyinput166, keyinput167, keyinput168, keyinput169;
  input keyinput170, keyinput171, keyinput172, keyinput173, keyinput174;
  input keyinput175, keyinput176, keyinput177, keyinput178, keyinput179;
  input keyinput180, keyinput181, keyinput182, keyinput183, keyinput184;
  input keyinput185, keyinput186, keyinput187, keyinput188, keyinput189;
  input keyinput190, keyinput191, keyinput192, keyinput193, keyinput194;
  input keyinput195, keyinput196, keyinput197, keyinput198, keyinput199;
  input keyinput200, keyinput201, keyinput202, keyinput203, keyinput204;
  input keyinput205, keyinput206, keyinput207, keyinput208, keyinput209;
  input keyinput210, keyinput211, keyinput212, keyinput213, keyinput214;
  input keyinput215, keyinput216, keyinput217, keyinput218, keyinput219;
  input keyinput220, keyinput221, keyinput222, keyinput223, keyinput224;
  input keyinput225, keyinput226, keyinput227, keyinput228, keyinput229;
  input keyinput230, keyinput231, keyinput232, keyinput233, keyinput234;
  input keyinput235, keyinput236, keyinput237, keyinput238, keyinput239;
  input keyinput240, keyinput241, keyinput242, keyinput243, keyinput244;
  input keyinput245, keyinput246, keyinput247, keyinput248, keyinput249;
  input keyinput250, keyinput251, keyinput252, keyinput253, keyinput254;
  input keyinput255;

  wire [0:255] keyinput_Wire_0;
  wire [0:123] KeyNOTWire_0;

input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;

output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;

wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877;

  nand NAND4_1 (keyinput_Wire_0[0], N1, N8, N13, N17);
  xor keyGate_0_0(KeyNOTWire_0[0], keyinput0, keyinput_Wire_0[0]);
  not KeyNOTGate_0_0(N269, KeyNOTWire_0[0]);
  nand NAND4_2 (keyinput_Wire_0[1], N1, N26, N13, N17);
  xnor keyGate_0_1(KeyNOTWire_0[1], keyinput1, keyinput_Wire_0[1]);
  not KeyNOTGate_0_1(N270, KeyNOTWire_0[1]);
  and AND3_3 (keyinput_Wire_0[2], N29, N36, N42);
  xor keyGate_0_2(KeyNOTWire_0[2], keyinput2, keyinput_Wire_0[2]);
  not KeyNOTGate_0_2(N273, KeyNOTWire_0[2]);
  and AND3_4 (keyinput_Wire_0[3], N1, N26, N51);
  xor keyGate_0_3(N276, keyinput3, keyinput_Wire_0[3]);
  nand NAND4_5 (keyinput_Wire_0[4], N1, N8, N51, N17);
  xor keyGate_0_4(N279, keyinput4, keyinput_Wire_0[4]);
  nand NAND4_6 (keyinput_Wire_0[5], N1, N8, N13, N55);
  xor keyGate_0_5(KeyNOTWire_0[3], keyinput5, keyinput_Wire_0[5]);
  not KeyNOTGate_0_3(N280, KeyNOTWire_0[3]);
  nand NAND4_7 (keyinput_Wire_0[6], N59, N42, N68, N72);
  xnor keyGate_0_6(KeyNOTWire_0[4], keyinput6, keyinput_Wire_0[6]);
  not KeyNOTGate_0_4(N284, KeyNOTWire_0[4]);
nand NAND2_8 (N285, N29, N68);
  nand NAND3_9 (keyinput_Wire_0[7], N59, N68, N74);
  xor keyGate_0_7(KeyNOTWire_0[5], keyinput7, keyinput_Wire_0[7]);
  not KeyNOTGate_0_5(N286, KeyNOTWire_0[5]);
and AND3_10 (N287, N29, N75, N80);
and AND3_11 (N290, N29, N75, N42);
  and AND3_12 (keyinput_Wire_0[8], N29, N36, N80);
  xor keyGate_0_8(N291, keyinput8, keyinput_Wire_0[8]);
  and AND3_13 (keyinput_Wire_0[9], N29, N36, N42);
  xor keyGate_0_9(N292, keyinput9, keyinput_Wire_0[9]);
  and AND3_14 (keyinput_Wire_0[10], N59, N75, N80);
  xor keyGate_0_10(KeyNOTWire_0[6], keyinput10, keyinput_Wire_0[10]);
  not KeyNOTGate_0_6(N293, KeyNOTWire_0[6]);
and AND3_15 (N294, N59, N75, N42);
  and AND3_16 (keyinput_Wire_0[11], N59, N36, N80);
  xnor keyGate_0_11(N295, keyinput11, keyinput_Wire_0[11]);
and AND3_17 (N296, N59, N36, N42);
  and AND2_18 (keyinput_Wire_0[12], N85, N86);
  xor keyGate_0_12(N297, keyinput12, keyinput_Wire_0[12]);
  or OR2_19 (keyinput_Wire_0[13], N87, N88);
  xor keyGate_0_13(KeyNOTWire_0[7], keyinput13, keyinput_Wire_0[13]);
  not KeyNOTGate_0_7(N298, KeyNOTWire_0[7]);
  nand NAND2_20 (keyinput_Wire_0[14], N91, N96);
  xor keyGate_0_14(KeyNOTWire_0[8], keyinput14, keyinput_Wire_0[14]);
  not KeyNOTGate_0_8(N301, KeyNOTWire_0[8]);
or OR2_21 (N302, N91, N96);
  nand NAND2_22 (keyinput_Wire_0[15], N101, N106);
  xor keyGate_0_15(N303, keyinput15, keyinput_Wire_0[15]);
or OR2_23 (N304, N101, N106);
nand NAND2_24 (N305, N111, N116);
  or OR2_25 (keyinput_Wire_0[16], N111, N116);
  xor keyGate_0_16(N306, keyinput16, keyinput_Wire_0[16]);
nand NAND2_26 (N307, N121, N126);
  or OR2_27 (keyinput_Wire_0[17], N121, N126);
  xnor keyGate_0_17(N308, keyinput17, keyinput_Wire_0[17]);
  and AND2_28 (keyinput_Wire_0[18], N8, N138);
  xnor keyGate_0_18(N309, keyinput18, keyinput_Wire_0[18]);
  not NOT1_29 (keyinput_Wire_0[19], N268);
  xnor keyGate_0_19(KeyNOTWire_0[9], keyinput19, keyinput_Wire_0[19]);
  not KeyNOTGate_0_9(N310, KeyNOTWire_0[9]);
and AND2_30 (N316, N51, N138);
  and AND2_31 (keyinput_Wire_0[20], N17, N138);
  xor keyGate_0_20(KeyNOTWire_0[10], keyinput20, keyinput_Wire_0[20]);
  not KeyNOTGate_0_10(N317, KeyNOTWire_0[10]);
and AND2_32 (N318, N152, N138);
  nand NAND2_33 (keyinput_Wire_0[21], N59, N156);
  xor keyGate_0_21(N319, keyinput21, keyinput_Wire_0[21]);
nor NOR2_34 (N322, N17, N42);
  and AND2_35 (keyinput_Wire_0[22], N17, N42);
  xnor keyGate_0_22(N323, keyinput22, keyinput_Wire_0[22]);
  nand NAND2_36 (keyinput_Wire_0[23], N159, N165);
  xnor keyGate_0_23(KeyNOTWire_0[11], keyinput23, keyinput_Wire_0[23]);
  not KeyNOTGate_0_11(N324, KeyNOTWire_0[11]);
  or OR2_37 (keyinput_Wire_0[24], N159, N165);
  xnor keyGate_0_24(N325, keyinput24, keyinput_Wire_0[24]);
  nand NAND2_38 (keyinput_Wire_0[25], N171, N177);
  xor keyGate_0_25(KeyNOTWire_0[12], keyinput25, keyinput_Wire_0[25]);
  not KeyNOTGate_0_12(N326, KeyNOTWire_0[12]);
  or OR2_39 (keyinput_Wire_0[26], N171, N177);
  xnor keyGate_0_26(N327, keyinput26, keyinput_Wire_0[26]);
  nand NAND2_40 (keyinput_Wire_0[27], N183, N189);
  xor keyGate_0_27(N328, keyinput27, keyinput_Wire_0[27]);
or OR2_41 (N329, N183, N189);
  nand NAND2_42 (keyinput_Wire_0[28], N195, N201);
  xnor keyGate_0_28(N330, keyinput28, keyinput_Wire_0[28]);
  or OR2_43 (keyinput_Wire_0[29], N195, N201);
  xor keyGate_0_29(N331, keyinput29, keyinput_Wire_0[29]);
  and AND2_44 (keyinput_Wire_0[30], N210, N91);
  xnor keyGate_0_30(N332, keyinput30, keyinput_Wire_0[30]);
  and AND2_45 (keyinput_Wire_0[31], N210, N96);
  xnor keyGate_0_31(KeyNOTWire_0[13], keyinput31, keyinput_Wire_0[31]);
  not KeyNOTGate_0_13(N333, KeyNOTWire_0[13]);
  and AND2_46 (keyinput_Wire_0[32], N210, N101);
  xor keyGate_0_32(N334, keyinput32, keyinput_Wire_0[32]);
  and AND2_47 (keyinput_Wire_0[33], N210, N106);
  xor keyGate_0_33(KeyNOTWire_0[14], keyinput33, keyinput_Wire_0[33]);
  not KeyNOTGate_0_14(N335, KeyNOTWire_0[14]);
  and AND2_48 (keyinput_Wire_0[34], N210, N111);
  xnor keyGate_0_34(N336, keyinput34, keyinput_Wire_0[34]);
  and AND2_49 (keyinput_Wire_0[35], N255, N259);
  xor keyGate_0_35(KeyNOTWire_0[15], keyinput35, keyinput_Wire_0[35]);
  not KeyNOTGate_0_15(N337, KeyNOTWire_0[15]);
  and AND2_50 (keyinput_Wire_0[36], N210, N116);
  xnor keyGate_0_36(N338, keyinput36, keyinput_Wire_0[36]);
and AND2_51 (N339, N255, N260);
and AND2_52 (N340, N210, N121);
and AND2_53 (N341, N255, N267);
  not NOT1_54 (keyinput_Wire_0[37], N269);
  xnor keyGate_0_37(KeyNOTWire_0[16], keyinput37, keyinput_Wire_0[37]);
  not KeyNOTGate_0_16(N342, KeyNOTWire_0[16]);
not NOT1_55 (N343, N273);
or OR2_56 (N344, N270, N273);
  not NOT1_57 (keyinput_Wire_0[38], N276);
  xor keyGate_0_38(N345, keyinput38, keyinput_Wire_0[38]);
  not NOT1_58 (keyinput_Wire_0[39], N276);
  xor keyGate_0_39(KeyNOTWire_0[17], keyinput39, keyinput_Wire_0[39]);
  not KeyNOTGate_0_17(N346, KeyNOTWire_0[17]);
  not NOT1_59 (keyinput_Wire_0[40], N279);
  xor keyGate_0_40(N347, keyinput40, keyinput_Wire_0[40]);
  nor NOR2_60 (keyinput_Wire_0[41], N280, N284);
  xor keyGate_0_41(KeyNOTWire_0[18], keyinput41, keyinput_Wire_0[41]);
  not KeyNOTGate_0_18(N348, KeyNOTWire_0[18]);
  or OR2_61 (keyinput_Wire_0[42], N280, N285);
  xor keyGate_0_42(N349, keyinput42, keyinput_Wire_0[42]);
or OR2_62 (N350, N280, N286);
  not NOT1_63 (keyinput_Wire_0[43], N293);
  xor keyGate_0_43(N351, keyinput43, keyinput_Wire_0[43]);
  not NOT1_64 (keyinput_Wire_0[44], N294);
  xor keyGate_0_44(KeyNOTWire_0[19], keyinput44, keyinput_Wire_0[44]);
  not KeyNOTGate_0_19(N352, KeyNOTWire_0[19]);
not NOT1_65 (N353, N295);
  not NOT1_66 (keyinput_Wire_0[45], N296);
  xor keyGate_0_45(KeyNOTWire_0[20], keyinput45, keyinput_Wire_0[45]);
  not KeyNOTGate_0_20(N354, KeyNOTWire_0[20]);
  nand NAND2_67 (keyinput_Wire_0[46], N89, N298);
  xor keyGate_0_46(N355, keyinput46, keyinput_Wire_0[46]);
  and AND2_68 (keyinput_Wire_0[47], N90, N298);
  xor keyGate_0_47(KeyNOTWire_0[21], keyinput47, keyinput_Wire_0[47]);
  not KeyNOTGate_0_21(N356, KeyNOTWire_0[21]);
nand NAND2_69 (N357, N301, N302);
nand NAND2_70 (N360, N303, N304);
  nand NAND2_71 (keyinput_Wire_0[48], N305, N306);
  xor keyGate_0_48(N363, keyinput48, keyinput_Wire_0[48]);
  nand NAND2_72 (keyinput_Wire_0[49], N307, N308);
  xor keyGate_0_49(KeyNOTWire_0[22], keyinput49, keyinput_Wire_0[49]);
  not KeyNOTGate_0_22(N366, KeyNOTWire_0[22]);
  not NOT1_73 (keyinput_Wire_0[50], N310);
  xor keyGate_0_50(N369, keyinput50, keyinput_Wire_0[50]);
  nor NOR2_74 (keyinput_Wire_0[51], N322, N323);
  xnor keyGate_0_51(N375, keyinput51, keyinput_Wire_0[51]);
  nand NAND2_75 (keyinput_Wire_0[52], N324, N325);
  xor keyGate_0_52(KeyNOTWire_0[23], keyinput52, keyinput_Wire_0[52]);
  not KeyNOTGate_0_23(N376, KeyNOTWire_0[23]);
  nand NAND2_76 (keyinput_Wire_0[53], N326, N327);
  xnor keyGate_0_53(N379, keyinput53, keyinput_Wire_0[53]);
  nand NAND2_77 (keyinput_Wire_0[54], N328, N329);
  xnor keyGate_0_54(KeyNOTWire_0[24], keyinput54, keyinput_Wire_0[54]);
  not KeyNOTGate_0_24(N382, KeyNOTWire_0[24]);
  nand NAND2_78 (keyinput_Wire_0[55], N330, N331);
  xnor keyGate_0_55(N385, keyinput55, keyinput_Wire_0[55]);
buf BUFF1_79 (N388, N290);
buf BUFF1_80 (KeyWire_0_1, N291);
  xor flip_it (N389, KeyWire_0_1, KeyWire_0_2 );
buf BUFF1_81 (N390, N292);
  buf BUFF1_82 (keyinput_Wire_1, N297);
  xor keyGate_1_1(N391, KeyWire_0_2, keyinput_Wire_1);
  or OR2_83 (keyinput_Wire_0[56], N270, N343);
  xor keyGate_0_56(KeyNOTWire_0[25], keyinput56, keyinput_Wire_0[56]);
  not KeyNOTGate_0_25(N392, KeyNOTWire_0[25]);
  not NOT1_84 (keyinput_Wire_0[57], N345);
  xor keyGate_0_57(KeyNOTWire_0[26], keyinput57, keyinput_Wire_0[57]);
  not KeyNOTGate_0_26(N393, KeyNOTWire_0[26]);
  not NOT1_85 (keyinput_Wire_0[58], N346);
  xor keyGate_0_58(KeyNOTWire_0[27], keyinput58, keyinput_Wire_0[58]);
  not KeyNOTGate_0_27(N399, KeyNOTWire_0[27]);
and AND2_86 (N400, N348, N73);
  not NOT1_87 (keyinput_Wire_0[59], N349);
  xor keyGate_0_59(KeyNOTWire_0[28], keyinput59, keyinput_Wire_0[59]);
  not KeyNOTGate_0_28(N401, KeyNOTWire_0[28]);
  not NOT1_88 (keyinput_Wire_0[60], N350);
  xnor keyGate_0_60(N402, keyinput60, keyinput_Wire_0[60]);
not NOT1_89 (N403, N355);
not NOT1_90 (N404, N357);
not NOT1_91 (N405, N360);
  and AND2_92 (keyinput_Wire_0[61], N357, N360);
  xnor keyGate_0_61(N406, keyinput61, keyinput_Wire_0[61]);
  not NOT1_93 (keyinput_Wire_0[62], N363);
  xor keyGate_0_62(N407, keyinput62, keyinput_Wire_0[62]);
  not NOT1_94 (keyinput_Wire_0[63], N366);
  xnor keyGate_0_63(KeyNOTWire_0[29], keyinput63, keyinput_Wire_0[63]);
  not KeyNOTGate_0_29(N408, KeyNOTWire_0[29]);
  and AND2_95 (keyinput_Wire_0[64], N363, N366);
  xor keyGate_0_64(N409, keyinput64, keyinput_Wire_0[64]);
  nand NAND2_96 (keyinput_Wire_0[65], N347, N352);
  xnor keyGate_0_65(N410, keyinput65, keyinput_Wire_0[65]);
  not NOT1_97 (keyinput_Wire_0[66], N376);
  xnor keyGate_0_66(KeyNOTWire_0[30], keyinput66, keyinput_Wire_0[66]);
  not KeyNOTGate_0_30(N411, KeyNOTWire_0[30]);
  not NOT1_98 (keyinput_Wire_0[67], N379);
  xor keyGate_0_67(KeyNOTWire_0[31], keyinput67, keyinput_Wire_0[67]);
  not KeyNOTGate_0_31(N412, KeyNOTWire_0[31]);
and AND2_99 (N413, N376, N379);
not NOT1_100 (N414, N382);
  not NOT1_101 (keyinput_Wire_0[68], N385);
  xnor keyGate_0_68(KeyNOTWire_0[32], keyinput68, keyinput_Wire_0[68]);
  not KeyNOTGate_0_32(N415, KeyNOTWire_0[32]);
and AND2_102 (N416, N382, N385);
  and AND2_103 (keyinput_Wire_0[69], N210, N369);
  xor keyGate_0_69(KeyNOTWire_0[33], keyinput69, keyinput_Wire_0[69]);
  not KeyNOTGate_0_33(N417, KeyNOTWire_0[33]);
buf BUFF1_104 (N418, N342);
buf BUFF1_105 (N419, N344);
buf BUFF1_106 (N420, N351);
buf BUFF1_107 (N421, N353);
buf BUFF1_108 (N422, N354);
buf BUFF1_109 (N423, N356);
not NOT1_110 (N424, N400);
  and AND2_111 (keyinput_Wire_0[70], N404, N405);
  xnor keyGate_0_70(KeyNOTWire_0[34], keyinput70, keyinput_Wire_0[70]);
  not KeyNOTGate_0_34(N425, KeyNOTWire_0[34]);
  and AND2_112 (keyinput_Wire_0[71], N407, N408);
  xnor keyGate_0_71(KeyNOTWire_0[35], keyinput71, keyinput_Wire_0[71]);
  not KeyNOTGate_0_35(N426, KeyNOTWire_0[35]);
  and AND3_113 (keyinput_Wire_0[72], N319, N393, N55);
  xor keyGate_0_72(KeyNOTWire_0[36], keyinput72, keyinput_Wire_0[72]);
  not KeyNOTGate_0_36(N427, KeyNOTWire_0[36]);
  and AND3_114 (keyinput_Wire_0[73], N393, N17, N287);
  xor keyGate_0_73(KeyNOTWire_0[37], keyinput73, keyinput_Wire_0[73]);
  not KeyNOTGate_0_37(N432, KeyNOTWire_0[37]);
  nand NAND3_115 (keyinput_Wire_0[74], N393, N287, N55);
  xnor keyGate_0_74(N437, keyinput74, keyinput_Wire_0[74]);
  nand NAND4_116 (keyinput_Wire_0[75], N375, N59, N156, N393);
  xor keyGate_0_75(KeyNOTWire_0[38], keyinput75, keyinput_Wire_0[75]);
  not KeyNOTGate_0_38(N442, KeyNOTWire_0[38]);
nand NAND3_117 (N443, N393, N319, N17);
  and AND2_118 (keyinput_Wire_0[76], N411, N412);
  xor keyGate_0_76(N444, keyinput76, keyinput_Wire_0[76]);
and AND2_119 (N445, N414, N415);
buf BUFF1_120 (N446, N392);
buf BUFF1_121 (N447, N399);
buf BUFF1_122 (N448, N401);
buf BUFF1_123 (N449, N402);
buf BUFF1_124 (N450, N403);
  not NOT1_125 (keyinput_Wire_0[77], N424);
  xnor keyGate_0_77(N451, keyinput77, keyinput_Wire_0[77]);
nor NOR2_126 (N460, N406, N425);
  nor NOR2_127 (keyinput_Wire_0[78], N409, N426);
  xor keyGate_0_78(N463, keyinput78, keyinput_Wire_0[78]);
  nand NAND2_128 (keyinput_Wire_0[79], N442, N410);
  xor keyGate_0_79(KeyNOTWire_0[39], keyinput79, keyinput_Wire_0[79]);
  not KeyNOTGate_0_39(N466, KeyNOTWire_0[39]);
and AND2_129 (N475, N143, N427);
  and AND2_130 (keyinput_Wire_0[80], N310, N432);
  xnor keyGate_0_80(KeyNOTWire_0[40], keyinput80, keyinput_Wire_0[80]);
  not KeyNOTGate_0_40(N476, KeyNOTWire_0[40]);
  and AND2_131 (keyinput_Wire_0[81], N146, N427);
  xnor keyGate_0_81(KeyNOTWire_0[41], keyinput81, keyinput_Wire_0[81]);
  not KeyNOTGate_0_41(N477, KeyNOTWire_0[41]);
  and AND2_132 (keyinput_Wire_0[82], N310, N432);
  xor keyGate_0_82(KeyNOTWire_0[42], keyinput82, keyinput_Wire_0[82]);
  not KeyNOTGate_0_42(N478, KeyNOTWire_0[42]);
  and AND2_133 (keyinput_Wire_0[83], N149, N427);
  xor keyGate_0_83(KeyNOTWire_0[43], keyinput83, keyinput_Wire_0[83]);
  not KeyNOTGate_0_43(N479, KeyNOTWire_0[43]);
and AND2_134 (N480, N310, N432);
  and AND2_135 (keyinput_Wire_0[84], N153, N427);
  xnor keyGate_0_84(KeyNOTWire_0[44], keyinput84, keyinput_Wire_0[84]);
  not KeyNOTGate_0_44(N481, KeyNOTWire_0[44]);
  and AND2_136 (keyinput_Wire_0[85], N310, N432);
  xor keyGate_0_85(N482, keyinput85, keyinput_Wire_0[85]);
nand NAND2_137 (N483, N443, N1);
  or OR2_138 (keyinput_Wire_0[86], N369, N437);
  xor keyGate_0_86(KeyNOTWire_0[45], keyinput86, keyinput_Wire_0[86]);
  not KeyNOTGate_0_45(N488, KeyNOTWire_0[45]);
  or OR2_139 (keyinput_Wire_0[87], N369, N437);
  xnor keyGate_0_87(N489, keyinput87, keyinput_Wire_0[87]);
  or OR2_140 (keyinput_Wire_0[88], N369, N437);
  xor keyGate_0_88(KeyNOTWire_0[46], keyinput88, keyinput_Wire_0[88]);
  not KeyNOTGate_0_46(N490, KeyNOTWire_0[46]);
  or OR2_141 (keyinput_Wire_0[89], N369, N437);
  xnor keyGate_0_89(KeyNOTWire_0[47], keyinput89, keyinput_Wire_0[89]);
  not KeyNOTGate_0_47(N491, KeyNOTWire_0[47]);
nor NOR2_142 (N492, N413, N444);
nor NOR2_143 (N495, N416, N445);
  nand NAND2_144 (keyinput_Wire_0[90], N130, N460);
  xnor keyGate_0_90(N498, keyinput90, keyinput_Wire_0[90]);
  or OR2_145 (keyinput_Wire_0[91], N130, N460);
  xor keyGate_0_91(KeyNOTWire_0[48], keyinput91, keyinput_Wire_0[91]);
  not KeyNOTGate_0_48(N499, KeyNOTWire_0[48]);
  nand NAND2_146 (keyinput_Wire_0[92], N463, N135);
  xor keyGate_0_92(N500, keyinput92, keyinput_Wire_0[92]);
  or OR2_147 (keyinput_Wire_0[93], N463, N135);
  xnor keyGate_0_93(KeyNOTWire_0[49], keyinput93, keyinput_Wire_0[93]);
  not KeyNOTGate_0_49(N501, KeyNOTWire_0[49]);
  and AND2_148 (keyinput_Wire_0[94], N91, N466);
  xor keyGate_0_94(N502, keyinput94, keyinput_Wire_0[94]);
  nor NOR2_149 (keyinput_Wire_0[95], N475, N476);
  xnor keyGate_0_95(KeyNOTWire_0[50], keyinput95, keyinput_Wire_0[95]);
  not KeyNOTGate_0_50(N503, KeyNOTWire_0[50]);
and AND2_150 (N504, N96, N466);
  nor NOR2_151 (keyinput_Wire_0[96], N477, N478);
  xor keyGate_0_96(KeyNOTWire_0[51], keyinput96, keyinput_Wire_0[96]);
  not KeyNOTGate_0_51(N505, KeyNOTWire_0[51]);
  and AND2_152 (keyinput_Wire_0[97], N101, N466);
  xnor keyGate_0_97(KeyNOTWire_0[52], keyinput97, keyinput_Wire_0[97]);
  not KeyNOTGate_0_52(N506, KeyNOTWire_0[52]);
  nor NOR2_153 (keyinput_Wire_0[98], N479, N480);
  xnor keyGate_0_98(KeyNOTWire_0[53], keyinput98, keyinput_Wire_0[98]);
  not KeyNOTGate_0_53(N507, KeyNOTWire_0[53]);
  and AND2_154 (keyinput_Wire_0[99], N106, N466);
  xnor keyGate_0_99(N508, keyinput99, keyinput_Wire_0[99]);
  nor NOR2_155 (keyinput_Wire_0[100], N481, N482);
  xor keyGate_0_100(KeyNOTWire_0[54], keyinput100, keyinput_Wire_0[100]);
  not KeyNOTGate_0_54(N509, KeyNOTWire_0[54]);
  and AND2_156 (keyinput_Wire_0[101], N143, N483);
  xnor keyGate_0_101(N510, keyinput101, keyinput_Wire_0[101]);
  and AND2_157 (keyinput_Wire_0[102], N111, N466);
  xor keyGate_0_102(KeyNOTWire_0[55], keyinput102, keyinput_Wire_0[102]);
  not KeyNOTGate_0_55(N511, KeyNOTWire_0[55]);
  and AND2_158 (keyinput_Wire_0[103], N146, N483);
  xor keyGate_0_103(N512, keyinput103, keyinput_Wire_0[103]);
  and AND2_159 (keyinput_Wire_0[104], N116, N466);
  xor keyGate_0_104(KeyNOTWire_0[56], keyinput104, keyinput_Wire_0[104]);
  not KeyNOTGate_0_56(N513, KeyNOTWire_0[56]);
  and AND2_160 (keyinput_Wire_0[105], N149, N483);
  xor keyGate_0_105(KeyNOTWire_0[57], keyinput105, keyinput_Wire_0[105]);
  not KeyNOTGate_0_57(N514, KeyNOTWire_0[57]);
  and AND2_161 (keyinput_Wire_0[106], N121, N466);
  xnor keyGate_0_106(N515, keyinput106, keyinput_Wire_0[106]);
and AND2_162 (N516, N153, N483);
and AND2_163 (N517, N126, N466);
  nand NAND2_164 (keyinput_Wire_0[107], N130, N492);
  xnor keyGate_0_107(N518, keyinput107, keyinput_Wire_0[107]);
  or OR2_165 (keyinput_Wire_0[108], N130, N492);
  xor keyGate_0_108(KeyNOTWire_0[58], keyinput108, keyinput_Wire_0[108]);
  not KeyNOTGate_0_58(N519, KeyNOTWire_0[58]);
  nand NAND2_166 (keyinput_Wire_0[109], N495, N207);
  xor keyGate_0_109(KeyNOTWire_0[59], keyinput109, keyinput_Wire_0[109]);
  not KeyNOTGate_0_59(N520, KeyNOTWire_0[59]);
or OR2_167 (N521, N495, N207);
  and AND2_168 (keyinput_Wire_0[110], N451, N159);
  xor keyGate_0_110(KeyNOTWire_0[60], keyinput110, keyinput_Wire_0[110]);
  not KeyNOTGate_0_60(N522, KeyNOTWire_0[60]);
  and AND2_169 (keyinput_Wire_0[111], N451, N165);
  xor keyGate_0_111(N523, keyinput111, keyinput_Wire_0[111]);
and AND2_170 (N524, N451, N171);
  and AND2_171 (keyinput_Wire_0[112], N451, N177);
  xor keyGate_0_112(KeyNOTWire_0[61], keyinput112, keyinput_Wire_0[112]);
  not KeyNOTGate_0_61(N525, KeyNOTWire_0[61]);
  and AND2_172 (keyinput_Wire_0[113], N451, N183);
  xor keyGate_0_113(N526, keyinput113, keyinput_Wire_0[113]);
nand NAND2_173 (N527, N451, N189);
  nand NAND2_174 (keyinput_Wire_0[114], N451, N195);
  xor keyGate_0_114(N528, keyinput114, keyinput_Wire_0[114]);
  nand NAND2_175 (keyinput_Wire_0[115], N451, N201);
  xor keyGate_0_115(N529, keyinput115, keyinput_Wire_0[115]);
  nand NAND2_176 (keyinput_Wire_0[116], N498, N499);
  xnor keyGate_0_116(N530, keyinput116, keyinput_Wire_0[116]);
  nand NAND2_177 (keyinput_Wire_0[117], N500, N501);
  xnor keyGate_0_117(KeyNOTWire_0[62], keyinput117, keyinput_Wire_0[117]);
  not KeyNOTGate_0_62(N533, KeyNOTWire_0[62]);
nor NOR2_178 (N536, N309, N502);
nor NOR2_179 (N537, N316, N504);
  nor NOR2_180 (keyinput_Wire_0[118], N317, N506);
  xnor keyGate_0_118(N538, keyinput118, keyinput_Wire_0[118]);
  nor NOR2_181 (keyinput_Wire_0[119], N318, N508);
  xnor keyGate_0_119(N539, keyinput119, keyinput_Wire_0[119]);
  nor NOR2_182 (keyinput_Wire_0[120], N510, N511);
  xnor keyGate_0_120(N540, keyinput120, keyinput_Wire_0[120]);
  nor NOR2_183 (keyinput_Wire_0[121], N512, N513);
  xnor keyGate_0_121(KeyNOTWire_0[63], keyinput121, keyinput_Wire_0[121]);
  not KeyNOTGate_0_63(N541, KeyNOTWire_0[63]);
nor NOR2_184 (N542, N514, N515);
  nor NOR2_185 (keyinput_Wire_0[122], N516, N517);
  xnor keyGate_0_122(KeyNOTWire_0[64], keyinput122, keyinput_Wire_0[122]);
  not KeyNOTGate_0_64(N543, KeyNOTWire_0[64]);
  nand NAND2_186 (keyinput_Wire_0[123], N518, N519);
  xor keyGate_0_123(N544, keyinput123, keyinput_Wire_0[123]);
nand NAND2_187 (N547, N520, N521);
  not NOT1_188 (keyinput_Wire_0[124], N530);
  xnor keyGate_0_124(N550, keyinput124, keyinput_Wire_0[124]);
  not NOT1_189 (keyinput_Wire_0[125], N533);
  xnor keyGate_0_125(KeyNOTWire_0[65], keyinput125, keyinput_Wire_0[125]);
  not KeyNOTGate_0_65(N551, KeyNOTWire_0[65]);
  and AND2_190 (keyinput_Wire_0[126], N530, N533);
  xor keyGate_0_126(N552, keyinput126, keyinput_Wire_0[126]);
  nand NAND2_191 (keyinput_Wire_0[127], N536, N503);
  xor keyGate_0_127(KeyNOTWire_0[66], keyinput127, keyinput_Wire_0[127]);
  not KeyNOTGate_0_66(N553, KeyNOTWire_0[66]);
  nand NAND2_192 (keyinput_Wire_0[128], N537, N505);
  xnor keyGate_0_128(N557, keyinput128, keyinput_Wire_0[128]);
  nand NAND2_193 (keyinput_Wire_0[129], N538, N507);
  xnor keyGate_0_129(KeyNOTWire_0[67], keyinput129, keyinput_Wire_0[129]);
  not KeyNOTGate_0_67(N561, KeyNOTWire_0[67]);
  nand NAND2_194 (keyinput_Wire_0[130], N539, N509);
  xnor keyGate_0_130(N565, keyinput130, keyinput_Wire_0[130]);
nand NAND2_195 (N569, N488, N540);
nand NAND2_196 (N573, N489, N541);
  nand NAND2_197 (keyinput_Wire_0[131], N490, N542);
  xnor keyGate_0_131(KeyNOTWire_0[68], keyinput131, keyinput_Wire_0[131]);
  not KeyNOTGate_0_68(N577, KeyNOTWire_0[68]);
  nand NAND2_198 (keyinput_Wire_0[132], N491, N543);
  xor keyGate_0_132(N581, keyinput132, keyinput_Wire_0[132]);
  not NOT1_199 (keyinput_Wire_0[133], N544);
  xnor keyGate_0_133(KeyNOTWire_0[69], keyinput133, keyinput_Wire_0[133]);
  not KeyNOTGate_0_69(N585, KeyNOTWire_0[69]);
  not NOT1_200 (keyinput_Wire_0[134], N547);
  xnor keyGate_0_134(KeyNOTWire_0[70], keyinput134, keyinput_Wire_0[134]);
  not KeyNOTGate_0_70(N586, KeyNOTWire_0[70]);
  and AND2_201 (keyinput_Wire_0[135], N544, N547);
  xor keyGate_0_135(KeyNOTWire_0[71], keyinput135, keyinput_Wire_0[135]);
  not KeyNOTGate_0_71(N587, KeyNOTWire_0[71]);
  and AND2_202 (keyinput_Wire_0[136], N550, N551);
  xnor keyGate_0_136(KeyNOTWire_0[72], keyinput136, keyinput_Wire_0[136]);
  not KeyNOTGate_0_72(N588, KeyNOTWire_0[72]);
  and AND2_203 (keyinput_Wire_0[137], N585, N586);
  xnor keyGate_0_137(N589, keyinput137, keyinput_Wire_0[137]);
nand NAND2_204 (N590, N553, N159);
  or OR2_205 (keyinput_Wire_0[138], N553, N159);
  xnor keyGate_0_138(N593, keyinput138, keyinput_Wire_0[138]);
and AND2_206 (N596, N246, N553);
  nand NAND2_207 (keyinput_Wire_0[139], N557, N165);
  xnor keyGate_0_139(N597, keyinput139, keyinput_Wire_0[139]);
  or OR2_208 (keyinput_Wire_0[140], N557, N165);
  xor keyGate_0_140(KeyNOTWire_0[73], keyinput140, keyinput_Wire_0[140]);
  not KeyNOTGate_0_73(N600, KeyNOTWire_0[73]);
  and AND2_209 (keyinput_Wire_0[141], N246, N557);
  xnor keyGate_0_141(N605, keyinput141, keyinput_Wire_0[141]);
  nand NAND2_210 (keyinput_Wire_0[142], N561, N171);
  xor keyGate_0_142(N606, keyinput142, keyinput_Wire_0[142]);
  or OR2_211 (keyinput_Wire_0[143], N561, N171);
  xnor keyGate_0_143(KeyNOTWire_0[74], keyinput143, keyinput_Wire_0[143]);
  not KeyNOTGate_0_74(N609, KeyNOTWire_0[74]);
  and AND2_212 (keyinput_Wire_0[144], N246, N561);
  xnor keyGate_0_144(N615, keyinput144, keyinput_Wire_0[144]);
nand NAND2_213 (N616, N565, N177);
or OR2_214 (N619, N565, N177);
  and AND2_215 (keyinput_Wire_0[145], N246, N565);
  xor keyGate_0_145(N624, keyinput145, keyinput_Wire_0[145]);
  nand NAND2_216 (keyinput_Wire_0[146], N569, N183);
  xor keyGate_0_146(KeyNOTWire_0[75], keyinput146, keyinput_Wire_0[146]);
  not KeyNOTGate_0_75(N625, KeyNOTWire_0[75]);
  or OR2_217 (keyinput_Wire_0[147], N569, N183);
  xnor keyGate_0_147(KeyNOTWire_0[76], keyinput147, keyinput_Wire_0[147]);
  not KeyNOTGate_0_76(N628, KeyNOTWire_0[76]);
  and AND2_218 (keyinput_Wire_0[148], N246, N569);
  xnor keyGate_0_148(N631, keyinput148, keyinput_Wire_0[148]);
nand NAND2_219 (N632, N573, N189);
  or OR2_220 (keyinput_Wire_0[149], N573, N189);
  xor keyGate_0_149(N635, keyinput149, keyinput_Wire_0[149]);
  and AND2_221 (keyinput_Wire_0[150], N246, N573);
  xor keyGate_0_150(N640, keyinput150, keyinput_Wire_0[150]);
  nand NAND2_222 (keyinput_Wire_0[151], N577, N195);
  xor keyGate_0_151(KeyNOTWire_0[77], keyinput151, keyinput_Wire_0[151]);
  not KeyNOTGate_0_77(N641, KeyNOTWire_0[77]);
  or OR2_223 (keyinput_Wire_0[152], N577, N195);
  xor keyGate_0_152(N644, keyinput152, keyinput_Wire_0[152]);
and AND2_224 (N650, N246, N577);
nand NAND2_225 (N651, N581, N201);
  or OR2_226 (keyinput_Wire_0[153], N581, N201);
  xnor keyGate_0_153(N654, keyinput153, keyinput_Wire_0[153]);
  and AND2_227 (keyinput_Wire_0[154], N246, N581);
  xor keyGate_0_154(N659, keyinput154, keyinput_Wire_0[154]);
  nor NOR2_228 (keyinput_Wire_0[155], N552, N588);
  xor keyGate_0_155(KeyNOTWire_0[78], keyinput155, keyinput_Wire_0[155]);
  not KeyNOTGate_0_78(N660, KeyNOTWire_0[78]);
nor NOR2_229 (N661, N587, N589);
  not NOT1_230 (keyinput_Wire_0[156], N590);
  xnor keyGate_0_156(N662, keyinput156, keyinput_Wire_0[156]);
  and AND2_231 (keyinput_Wire_0[157], N593, N590);
  xor keyGate_0_157(N665, keyinput157, keyinput_Wire_0[157]);
nor NOR2_232 (N669, N596, N522);
  not NOT1_233 (keyinput_Wire_0[158], N597);
  xnor keyGate_0_158(N670, keyinput158, keyinput_Wire_0[158]);
  and AND2_234 (keyinput_Wire_0[159], N600, N597);
  xor keyGate_0_159(N673, keyinput159, keyinput_Wire_0[159]);
  nor NOR2_235 (keyinput_Wire_0[160], N605, N523);
  xnor keyGate_0_160(KeyNOTWire_0[79], keyinput160, keyinput_Wire_0[160]);
  not KeyNOTGate_0_79(N677, KeyNOTWire_0[79]);
  not NOT1_236 (keyinput_Wire_0[161], N606);
  xnor keyGate_0_161(KeyNOTWire_0[80], keyinput161, keyinput_Wire_0[161]);
  not KeyNOTGate_0_80(N678, KeyNOTWire_0[80]);
  and AND2_237 (keyinput_Wire_0[162], N609, N606);
  xnor keyGate_0_162(KeyNOTWire_0[81], keyinput162, keyinput_Wire_0[162]);
  not KeyNOTGate_0_81(N682, KeyNOTWire_0[81]);
  nor NOR2_238 (keyinput_Wire_0[163], N615, N524);
  xnor keyGate_0_163(KeyNOTWire_0[82], keyinput163, keyinput_Wire_0[163]);
  not KeyNOTGate_0_82(N686, KeyNOTWire_0[82]);
  not NOT1_239 (keyinput_Wire_0[164], N616);
  xnor keyGate_0_164(N687, keyinput164, keyinput_Wire_0[164]);
  and AND2_240 (keyinput_Wire_0[165], N619, N616);
  xor keyGate_0_165(KeyNOTWire_0[83], keyinput165, keyinput_Wire_0[165]);
  not KeyNOTGate_0_83(N692, KeyNOTWire_0[83]);
  nor NOR2_241 (keyinput_Wire_0[166], N624, N525);
  xnor keyGate_0_166(KeyNOTWire_0[84], keyinput166, keyinput_Wire_0[166]);
  not KeyNOTGate_0_84(N696, KeyNOTWire_0[84]);
  not NOT1_242 (keyinput_Wire_0[167], N625);
  xnor keyGate_0_167(N697, keyinput167, keyinput_Wire_0[167]);
  and AND2_243 (keyinput_Wire_0[168], N628, N625);
  xor keyGate_0_168(N700, keyinput168, keyinput_Wire_0[168]);
  nor NOR2_244 (keyinput_Wire_0[169], N631, N526);
  xor keyGate_0_169(N704, keyinput169, keyinput_Wire_0[169]);
not NOT1_245 (N705, N632);
  and AND2_246 (keyinput_Wire_0[170], N635, N632);
  xor keyGate_0_170(KeyNOTWire_0[85], keyinput170, keyinput_Wire_0[170]);
  not KeyNOTGate_0_85(N708, KeyNOTWire_0[85]);
  nor NOR2_247 (keyinput_Wire_0[171], N337, N640);
  xnor keyGate_0_171(KeyNOTWire_0[86], keyinput171, keyinput_Wire_0[171]);
  not KeyNOTGate_0_86(N712, KeyNOTWire_0[86]);
  not NOT1_248 (keyinput_Wire_0[172], N641);
  xnor keyGate_0_172(KeyNOTWire_0[87], keyinput172, keyinput_Wire_0[172]);
  not KeyNOTGate_0_87(N713, KeyNOTWire_0[87]);
and AND2_249 (N717, N644, N641);
  nor NOR2_250 (keyinput_Wire_0[173], N339, N650);
  xnor keyGate_0_173(KeyNOTWire_0[88], keyinput173, keyinput_Wire_0[173]);
  not KeyNOTGate_0_88(N721, KeyNOTWire_0[88]);
not NOT1_251 (N722, N651);
  and AND2_252 (keyinput_Wire_0[174], N654, N651);
  xor keyGate_0_174(KeyNOTWire_0[89], keyinput174, keyinput_Wire_0[174]);
  not KeyNOTGate_0_89(N727, KeyNOTWire_0[89]);
  nor NOR2_253 (keyinput_Wire_0[175], N341, N659);
  xnor keyGate_0_175(N731, keyinput175, keyinput_Wire_0[175]);
  nand NAND2_254 (keyinput_Wire_0[176], N654, N261);
  xnor keyGate_0_176(N732, keyinput176, keyinput_Wire_0[176]);
  nand NAND3_255 (keyinput_Wire_0[177], N644, N654, N261);
  xor keyGate_0_177(N733, keyinput177, keyinput_Wire_0[177]);
  nand NAND4_256 (keyinput_Wire_0[178], N635, N644, N654, N261);
  xnor keyGate_0_178(KeyNOTWire_0[90], keyinput178, keyinput_Wire_0[178]);
  not KeyNOTGate_0_90(N734, KeyNOTWire_0[90]);
not NOT1_257 (N735, N662);
and AND2_258 (N736, N228, N665);
  and AND2_259 (keyinput_Wire_0[179], N237, N662);
  xnor keyGate_0_179(N737, keyinput179, keyinput_Wire_0[179]);
not NOT1_260 (N738, N670);
  and AND2_261 (keyinput_Wire_0[180], N228, N673);
  xnor keyGate_0_180(N739, keyinput180, keyinput_Wire_0[180]);
  and AND2_262 (keyinput_Wire_0[181], N237, N670);
  xor keyGate_0_181(N740, keyinput181, keyinput_Wire_0[181]);
  not NOT1_263 (keyinput_Wire_0[182], N678);
  xor keyGate_0_182(KeyNOTWire_0[91], keyinput182, keyinput_Wire_0[182]);
  not KeyNOTGate_0_91(N741, KeyNOTWire_0[91]);
  and AND2_264 (keyinput_Wire_0[183], N228, N682);
  xor keyGate_0_183(N742, keyinput183, keyinput_Wire_0[183]);
and AND2_265 (N743, N237, N678);
  not NOT1_266 (keyinput_Wire_0[184], N687);
  xor keyGate_0_184(N744, keyinput184, keyinput_Wire_0[184]);
and AND2_267 (N745, N228, N692);
and AND2_268 (N746, N237, N687);
  not NOT1_269 (keyinput_Wire_0[185], N697);
  xor keyGate_0_185(KeyNOTWire_0[92], keyinput185, keyinput_Wire_0[185]);
  not KeyNOTGate_0_92(N747, KeyNOTWire_0[92]);
  and AND2_270 (keyinput_Wire_0[186], N228, N700);
  xnor keyGate_0_186(KeyNOTWire_0[93], keyinput186, keyinput_Wire_0[186]);
  not KeyNOTGate_0_93(N748, KeyNOTWire_0[93]);
and AND2_271 (N749, N237, N697);
not NOT1_272 (N750, N705);
  and AND2_273 (keyinput_Wire_0[187], N228, N708);
  xnor keyGate_0_187(N751, keyinput187, keyinput_Wire_0[187]);
  and AND2_274 (keyinput_Wire_0[188], N237, N705);
  xnor keyGate_0_188(N752, keyinput188, keyinput_Wire_0[188]);
  not NOT1_275 (keyinput_Wire_0[189], N713);
  xor keyGate_0_189(N753, keyinput189, keyinput_Wire_0[189]);
  and AND2_276 (keyinput_Wire_0[190], N228, N717);
  xnor keyGate_0_190(N754, keyinput190, keyinput_Wire_0[190]);
and AND2_277 (N755, N237, N713);
not NOT1_278 (N756, N722);
  nor NOR2_279 (keyinput_Wire_0[191], N727, N261);
  xor keyGate_0_191(N757, keyinput191, keyinput_Wire_0[191]);
  and AND2_280 (keyinput_Wire_0[192], N727, N261);
  xor keyGate_0_192(N758, keyinput192, keyinput_Wire_0[192]);
and AND2_281 (N759, N228, N727);
  and AND2_282 (keyinput_Wire_0[193], N237, N722);
  xnor keyGate_0_193(KeyNOTWire_0[94], keyinput193, keyinput_Wire_0[193]);
  not KeyNOTGate_0_94(N760, KeyNOTWire_0[94]);
  nand NAND2_283 (keyinput_Wire_0[194], N644, N722);
  xor keyGate_0_194(KeyNOTWire_0[95], keyinput194, keyinput_Wire_0[194]);
  not KeyNOTGate_0_95(N761, KeyNOTWire_0[95]);
nand NAND2_284 (N762, N635, N713);
nand NAND3_285 (N763, N635, N644, N722);
  nand NAND2_286 (keyinput_Wire_0[195], N609, N687);
  xnor keyGate_0_195(N764, keyinput195, keyinput_Wire_0[195]);
nand NAND2_287 (N765, N600, N678);
  nand NAND3_288 (keyinput_Wire_0[196], N600, N609, N687);
  xnor keyGate_0_196(N766, keyinput196, keyinput_Wire_0[196]);
buf BUFF1_289 (N767, N660);
buf BUFF1_290 (N768, N661);
  nor NOR2_291 (keyinput_Wire_0[197], N736, N737);
  xor keyGate_0_197(N769, keyinput197, keyinput_Wire_0[197]);
nor NOR2_292 (N770, N739, N740);
  nor NOR2_293 (keyinput_Wire_0[198], N742, N743);
  xor keyGate_0_198(KeyNOTWire_0[96], keyinput198, keyinput_Wire_0[198]);
  not KeyNOTGate_0_96(N771, KeyNOTWire_0[96]);
nor NOR2_294 (N772, N745, N746);
nand NAND4_295 (N773, N750, N762, N763, N734);
  nor NOR2_296 (keyinput_Wire_0[199], N748, N749);
  xor keyGate_0_199(KeyNOTWire_0[97], keyinput199, keyinput_Wire_0[199]);
  not KeyNOTGate_0_97(N777, KeyNOTWire_0[97]);
  nand NAND3_297 (keyinput_Wire_0[200], N753, N761, N733);
  xor keyGate_0_200(KeyNOTWire_0[98], keyinput200, keyinput_Wire_0[200]);
  not KeyNOTGate_0_98(N778, KeyNOTWire_0[98]);
nor NOR2_298 (N781, N751, N752);
  nand NAND2_299 (keyinput_Wire_0[201], N756, N732);
  xor keyGate_0_201(N782, keyinput201, keyinput_Wire_0[201]);
  nor NOR2_300 (keyinput_Wire_0[202], N754, N755);
  xnor keyGate_0_202(KeyNOTWire_0[99], keyinput202, keyinput_Wire_0[202]);
  not KeyNOTGate_0_99(N785, KeyNOTWire_0[99]);
  nor NOR2_301 (keyinput_Wire_0[203], N757, N758);
  xor keyGate_0_203(KeyNOTWire_0[100], keyinput203, keyinput_Wire_0[203]);
  not KeyNOTGate_0_100(N786, KeyNOTWire_0[100]);
  nor NOR2_302 (keyinput_Wire_0[204], N759, N760);
  xnor keyGate_0_204(N787, keyinput204, keyinput_Wire_0[204]);
  nor NOR2_303 (keyinput_Wire_0[205], N700, N773);
  xnor keyGate_0_205(N788, keyinput205, keyinput_Wire_0[205]);
  and AND2_304 (keyinput_Wire_0[206], N700, N773);
  xor keyGate_0_206(KeyNOTWire_0[101], keyinput206, keyinput_Wire_0[206]);
  not KeyNOTGate_0_101(N789, KeyNOTWire_0[101]);
  nor NOR2_305 (keyinput_Wire_0[207], N708, N778);
  xnor keyGate_0_207(N790, keyinput207, keyinput_Wire_0[207]);
  and AND2_306 (keyinput_Wire_0[208], N708, N778);
  xor keyGate_0_208(KeyNOTWire_0[102], keyinput208, keyinput_Wire_0[208]);
  not KeyNOTGate_0_102(N791, KeyNOTWire_0[102]);
  nor NOR2_307 (keyinput_Wire_0[209], N717, N782);
  xnor keyGate_0_209(KeyNOTWire_0[103], keyinput209, keyinput_Wire_0[209]);
  not KeyNOTGate_0_103(N792, KeyNOTWire_0[103]);
  and AND2_308 (keyinput_Wire_0[210], N717, N782);
  xor keyGate_0_210(KeyNOTWire_0[104], keyinput210, keyinput_Wire_0[210]);
  not KeyNOTGate_0_104(N793, KeyNOTWire_0[104]);
  and AND2_309 (keyinput_Wire_0[211], N219, N786);
  xor keyGate_0_211(N794, keyinput211, keyinput_Wire_0[211]);
nand NAND2_310 (N795, N628, N773);
nand NAND2_311 (N796, N795, N747);
nor NOR2_312 (N802, N788, N789);
nor NOR2_313 (N803, N790, N791);
  nor NOR2_314 (keyinput_Wire_0[212], N792, N793);
  xnor keyGate_0_212(N804, keyinput212, keyinput_Wire_0[212]);
  nor NOR2_315 (keyinput_Wire_0[213], N340, N794);
  xnor keyGate_0_213(KeyNOTWire_0[105], keyinput213, keyinput_Wire_0[213]);
  not KeyNOTGate_0_105(N805, KeyNOTWire_0[105]);
nor NOR2_316 (N806, N692, N796);
  and AND2_317 (keyinput_Wire_0[214], N692, N796);
  xnor keyGate_0_214(KeyNOTWire_0[106], keyinput214, keyinput_Wire_0[214]);
  not KeyNOTGate_0_106(N807, KeyNOTWire_0[106]);
  and AND2_318 (keyinput_Wire_0[215], N219, N802);
  xnor keyGate_0_215(N808, keyinput215, keyinput_Wire_0[215]);
  and AND2_319 (keyinput_Wire_0[216], N219, N803);
  xor keyGate_0_216(KeyNOTWire_0[107], keyinput216, keyinput_Wire_0[216]);
  not KeyNOTGate_0_107(N809, KeyNOTWire_0[107]);
and AND2_320 (N810, N219, N804);
  nand NAND4_321 (keyinput_Wire_0[217], N805, N787, N731, N529);
  xnor keyGate_0_217(N811, keyinput217, keyinput_Wire_0[217]);
nand NAND2_322 (N812, N619, N796);
nand NAND3_323 (N813, N609, N619, N796);
  nand NAND4_324 (keyinput_Wire_0[218], N600, N609, N619, N796);
  xor keyGate_0_218(KeyNOTWire_0[108], keyinput218, keyinput_Wire_0[218]);
  not KeyNOTGate_0_108(N814, KeyNOTWire_0[108]);
  nand NAND4_325 (keyinput_Wire_0[219], N738, N765, N766, N814);
  xor keyGate_0_219(KeyNOTWire_0[109], keyinput219, keyinput_Wire_0[219]);
  not KeyNOTGate_0_109(N815, KeyNOTWire_0[109]);
  nand NAND3_326 (keyinput_Wire_0[220], N741, N764, N813);
  xnor keyGate_0_220(N819, keyinput220, keyinput_Wire_0[220]);
  nand NAND2_327 (keyinput_Wire_0[221], N744, N812);
  xnor keyGate_0_221(KeyNOTWire_0[110], keyinput221, keyinput_Wire_0[221]);
  not KeyNOTGate_0_110(N822, KeyNOTWire_0[110]);
  nor NOR2_328 (keyinput_Wire_0[222], N806, N807);
  xnor keyGate_0_222(KeyNOTWire_0[111], keyinput222, keyinput_Wire_0[222]);
  not KeyNOTGate_0_111(N825, KeyNOTWire_0[111]);
nor NOR2_329 (N826, N335, N808);
  nor NOR2_330 (keyinput_Wire_0[223], N336, N809);
  xor keyGate_0_223(N827, keyinput223, keyinput_Wire_0[223]);
  nor NOR2_331 (keyinput_Wire_0[224], N338, N810);
  xnor keyGate_0_224(KeyNOTWire_0[112], keyinput224, keyinput_Wire_0[224]);
  not KeyNOTGate_0_112(N828, KeyNOTWire_0[112]);
  not NOT1_332 (keyinput_Wire_0[225], N811);
  xor keyGate_0_225(KeyNOTWire_0[113], keyinput225, keyinput_Wire_0[225]);
  not KeyNOTGate_0_113(N829, KeyNOTWire_0[113]);
  nor NOR2_333 (keyinput_Wire_0[226], N665, N815);
  xnor keyGate_0_226(N830, keyinput226, keyinput_Wire_0[226]);
  and AND2_334 (keyinput_Wire_0[227], N665, N815);
  xor keyGate_0_227(N831, keyinput227, keyinput_Wire_0[227]);
  nor NOR2_335 (keyinput_Wire_0[228], N673, N819);
  xor keyGate_0_228(KeyNOTWire_0[114], keyinput228, keyinput_Wire_0[228]);
  not KeyNOTGate_0_114(N832, KeyNOTWire_0[114]);
  and AND2_336 (keyinput_Wire_0[229], N673, N819);
  xor keyGate_0_229(KeyNOTWire_0[115], keyinput229, keyinput_Wire_0[229]);
  not KeyNOTGate_0_115(N833, KeyNOTWire_0[115]);
nor NOR2_337 (N834, N682, N822);
and AND2_338 (N835, N682, N822);
and AND2_339 (N836, N219, N825);
nand NAND3_340 (N837, N826, N777, N704);
  nand NAND4_341 (keyinput_Wire_0[230], N827, N781, N712, N527);
  xnor keyGate_0_230(N838, keyinput230, keyinput_Wire_0[230]);
  nand NAND4_342 (keyinput_Wire_0[231], N828, N785, N721, N528);
  xor keyGate_0_231(N839, keyinput231, keyinput_Wire_0[231]);
  not NOT1_343 (keyinput_Wire_0[232], N829);
  xnor keyGate_0_232(N840, keyinput232, keyinput_Wire_0[232]);
  nand NAND2_344 (keyinput_Wire_0[233], N815, N593);
  xnor keyGate_0_233(KeyNOTWire_0[116], keyinput233, keyinput_Wire_0[233]);
  not KeyNOTGate_0_116(N841, KeyNOTWire_0[116]);
nor NOR2_345 (N842, N830, N831);
  nor NOR2_346 (keyinput_Wire_0[234], N832, N833);
  xor keyGate_0_234(N843, keyinput234, keyinput_Wire_0[234]);
  nor NOR2_347 (keyinput_Wire_0[235], N834, N835);
  xnor keyGate_0_235(KeyNOTWire_0[117], keyinput235, keyinput_Wire_0[235]);
  not KeyNOTGate_0_117(N844, KeyNOTWire_0[117]);
  nor NOR2_348 (keyinput_Wire_0[236], N334, N836);
  xnor keyGate_0_236(N845, keyinput236, keyinput_Wire_0[236]);
  not NOT1_349 (keyinput_Wire_0[237], N837);
  xor keyGate_0_237(N846, keyinput237, keyinput_Wire_0[237]);
not NOT1_350 (N847, N838);
not NOT1_351 (N848, N839);
and AND2_352 (N849, N735, N841);
buf BUFF1_353 (N850, N840);
  and AND2_354 (keyinput_Wire_0[238], N219, N842);
  xor keyGate_0_238(KeyNOTWire_0[118], keyinput238, keyinput_Wire_0[238]);
  not KeyNOTGate_0_118(N851, KeyNOTWire_0[118]);
  and AND2_355 (keyinput_Wire_0[239], N219, N843);
  xnor keyGate_0_239(N852, keyinput239, keyinput_Wire_0[239]);
  and AND2_356 (keyinput_Wire_0[240], N219, N844);
  xnor keyGate_0_240(KeyNOTWire_0[119], keyinput240, keyinput_Wire_0[240]);
  not KeyNOTGate_0_119(N853, KeyNOTWire_0[119]);
  nand NAND3_357 (keyinput_Wire_0[241], N845, N772, N696);
  xnor keyGate_0_241(N854, keyinput241, keyinput_Wire_0[241]);
  not NOT1_358 (keyinput_Wire_0[242], N846);
  xor keyGate_0_242(N855, keyinput242, keyinput_Wire_0[242]);
  not NOT1_359 (keyinput_Wire_0[243], N847);
  xor keyGate_0_243(KeyNOTWire_0[120], keyinput243, keyinput_Wire_0[243]);
  not KeyNOTGate_0_120(N856, KeyNOTWire_0[120]);
  not NOT1_360 (keyinput_Wire_0[244], N848);
  xor keyGate_0_244(KeyNOTWire_0[121], keyinput244, keyinput_Wire_0[244]);
  not KeyNOTGate_0_121(N857, KeyNOTWire_0[121]);
  not NOT1_361 (keyinput_Wire_0[245], N849);
  xnor keyGate_0_245(N858, keyinput245, keyinput_Wire_0[245]);
  nor NOR2_362 (keyinput_Wire_0[246], N417, N851);
  xnor keyGate_0_246(N859, keyinput246, keyinput_Wire_0[246]);
  nor NOR2_363 (keyinput_Wire_0[247], N332, N852);
  xnor keyGate_0_247(N860, keyinput247, keyinput_Wire_0[247]);
  nor NOR2_364 (keyinput_Wire_0[248], N333, N853);
  xnor keyGate_0_248(N861, keyinput248, keyinput_Wire_0[248]);
  not NOT1_365 (keyinput_Wire_0[249], N854);
  xor keyGate_0_249(N862, keyinput249, keyinput_Wire_0[249]);
buf BUFF1_366 (N863, N855);
buf BUFF1_367 (N864, N856);
buf BUFF1_368 (N865, N857);
buf BUFF1_369 (N866, N858);
nand NAND3_370 (N867, N859, N769, N669);
  nand NAND3_371 (keyinput_Wire_0[250], N860, N770, N677);
  xnor keyGate_0_250(N868, keyinput250, keyinput_Wire_0[250]);
nand NAND3_372 (N869, N861, N771, N686);
not NOT1_373 (N870, N862);
  not NOT1_374 (keyinput_Wire_0[251], N867);
  xor keyGate_0_251(N871, keyinput251, keyinput_Wire_0[251]);
  not NOT1_375 (keyinput_Wire_0[252], N868);
  xor keyGate_0_252(N872, keyinput252, keyinput_Wire_0[252]);
not NOT1_376 (N873, N869);
buf BUFF1_377 (N874, N870);
  not NOT1_378 (keyinput_Wire_0[253], N871);
  xnor keyGate_0_253(KeyNOTWire_0[122], keyinput253, keyinput_Wire_0[253]);
  not KeyNOTGate_0_122(N875, KeyNOTWire_0[122]);
  not NOT1_379 (keyinput_Wire_0[254], N872);
  xor keyGate_0_254(KeyNOTWire_0[123], keyinput254, keyinput_Wire_0[254]);
  not KeyNOTGate_0_123(N876, KeyNOTWire_0[123]);
  not NOT1_380 (keyinput_Wire_0[255], N873);
  xor keyGate_0_255(N877, keyinput255, keyinput_Wire_0[255]);
buf BUFF1_381 (N878, N875);
buf BUFF1_382 (N879, N876);
buf BUFF1_383 (N880, N877);

AntiSAT some_name( KeyWire_0_2, N26, N189, N138, N68, N143, N91, N159, N101, N219, N156, N116, N72, N90, N121, N246, N135, N86, N42, N130, N13, N195, N29, N106, N75, N87, N8, N85, N126, N51, N259, N152, N55, N171, N73, N165, N177, N201, N153, N1, N74, N80, N261, N237, N146, N96, N268, N59, N17, N89, N88, N111, N149, N36, N255, N267, N228, N207, N210, N183, N260, keyinput256, keyinput257, keyinput258, keyinput259, keyinput260, keyinput261, keyinput262, keyinput263, keyinput264, keyinput265, keyinput266, keyinput267, keyinput268, keyinput269, keyinput270, keyinput271, keyinput272, keyinput273, keyinput274, keyinput275, keyinput276, keyinput277, keyinput278, keyinput279, keyinput280, keyinput281, keyinput282, keyinput283, keyinput284, keyinput285, keyinput286, keyinput287, keyinput288, keyinput289, keyinput290, keyinput291, keyinput292, keyinput293, keyinput294, keyinput295, keyinput296, keyinput297, keyinput298, keyinput299, keyinput300, keyinput301, keyinput302, keyinput303, keyinput304, keyinput305, keyinput306, keyinput307, keyinput308, keyinput309, keyinput310, keyinput311, keyinput312, keyinput313, keyinput314, keyinput315, keyinput316, keyinput317, keyinput318, keyinput319, keyinput320, keyinput321, keyinput322, keyinput323, keyinput324, keyinput325, keyinput326, keyinput327, keyinput328, keyinput329, keyinput330, keyinput331, keyinput332, keyinput333, keyinput334, keyinput335, keyinput336, keyinput337, keyinput338, keyinput339, keyinput340, keyinput341, keyinput342, keyinput343, keyinput344, keyinput345, keyinput346, keyinput347, keyinput348, keyinput349, keyinput350, keyinput351, keyinput352, keyinput353, keyinput354, keyinput355, keyinput356, keyinput357, keyinput358, keyinput359, keyinput360, keyinput361, keyinput362, keyinput363, keyinput364, keyinput365, keyinput366, keyinput367, keyinput368, keyinput369, keyinput370, keyinput371, keyinput372, keyinput373, keyinput374, keyinput375,
       keyinput376, keyinput377, keyinput378, keyinput379, keyinput380,
       keyinput381, keyinput382, keyinput383, keyinput384, keyinput385,
       keyinput386, keyinput387, keyinput388, keyinput389, keyinput390,
       keyinput391, keyinput392, keyinput393, keyinput394, keyinput395,
       keyinput396, keyinput397, keyinput398, keyinput399, keyinput400,
       keyinput401, keyinput402, keyinput403, keyinput404, keyinput405,
       keyinput406, keyinput407, keyinput408, keyinput409, keyinput410,
       keyinput411, keyinput412, keyinput413, keyinput414, keyinput415,
       keyinput416, keyinput417, keyinput418, keyinput419, keyinput420,
       keyinput421, keyinput422, keyinput423, keyinput424, keyinput425,
       keyinput426, keyinput427, keyinput428, keyinput429, keyinput430,
       keyinput431, keyinput432, keyinput433, keyinput434, keyinput435);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N26, N189, N138, N68, N143, N91, N159, N101, N219, N156, N116, N72, N90, N121, N246, N135, N86, N42, N130, N13, N195, N29, N106, N75, N87, N8, N85, N126, N51, N259, N152, N55, N171, N73, N165, N177, N201, N153, N1, N74, N80, N261, N237, N146, N96, N268, N59, N17, N89, N88, N111, N149, N36, N255, N267, N228, N207, N210, N183, N260, keyinput256, keyinput257, keyinput258, keyinput259, keyinput260, keyinput261, keyinput262, keyinput263, keyinput264, keyinput265, keyinput266, keyinput267, keyinput268, keyinput269, keyinput270, keyinput271, keyinput272, keyinput273, keyinput274, keyinput275, keyinput276, keyinput277, keyinput278, keyinput279, keyinput280, keyinput281, keyinput282, keyinput283, keyinput284, keyinput285, keyinput286, keyinput287, keyinput288, keyinput289, keyinput290, keyinput291, keyinput292, keyinput293, keyinput294, keyinput295, keyinput296, keyinput297, keyinput298, keyinput299, keyinput300, keyinput301, keyinput302, keyinput303, keyinput304, keyinput305, keyinput306, keyinput307, keyinput308, keyinput309, keyinput310, keyinput311, keyinput312, keyinput313, keyinput314, keyinput315, keyinput316, keyinput317, keyinput318, keyinput319, keyinput320, keyinput321, keyinput322, keyinput323, keyinput324, keyinput325, keyinput326, keyinput327, keyinput328, keyinput329, keyinput330, keyinput331, keyinput332, keyinput333, keyinput334, keyinput335, keyinput336, keyinput337, keyinput338, keyinput339, keyinput340, keyinput341, keyinput342, keyinput343, keyinput344, keyinput345, keyinput346, keyinput347, keyinput348, keyinput349, keyinput350, keyinput351, keyinput352, keyinput353, keyinput354, keyinput355, keyinput356, keyinput357, keyinput358, keyinput359, keyinput360, keyinput361, keyinput362, keyinput363, keyinput364, keyinput365, keyinput366, keyinput367, keyinput368, keyinput369, keyinput370, keyinput371, keyinput372, keyinput373, keyinput374, keyinput375 ,
        keyinput376, keyinput377, keyinput378, keyinput379, keyinput380,
        keyinput381, keyinput382, keyinput383, keyinput384, keyinput385,
        keyinput386, keyinput387, keyinput388, keyinput389, keyinput390,
        keyinput391, keyinput392, keyinput393, keyinput394, keyinput395,
        keyinput396, keyinput397, keyinput398, keyinput399, keyinput400,
        keyinput401, keyinput402, keyinput403, keyinput404, keyinput405,
        keyinput406, keyinput407, keyinput408, keyinput409, keyinput410,
        keyinput411, keyinput412, keyinput413, keyinput414, keyinput415,
        keyinput416, keyinput417, keyinput418, keyinput419, keyinput420,
        keyinput421, keyinput422, keyinput423, keyinput424, keyinput425,
        keyinput426, keyinput427, keyinput428, keyinput429, keyinput430,
        keyinput431, keyinput432, keyinput433, keyinput434, keyinput435);

  input keyinput376, keyinput377, keyinput378, keyinput379, keyinput380;
  input keyinput381, keyinput382, keyinput383, keyinput384, keyinput385;
  input keyinput386, keyinput387, keyinput388, keyinput389, keyinput390;
  input keyinput391, keyinput392, keyinput393, keyinput394, keyinput395;
  input keyinput396, keyinput397, keyinput398, keyinput399, keyinput400;
  input keyinput401, keyinput402, keyinput403, keyinput404, keyinput405;
  input keyinput406, keyinput407, keyinput408, keyinput409, keyinput410;
  input keyinput411, keyinput412, keyinput413, keyinput414, keyinput415;
  input keyinput416, keyinput417, keyinput418, keyinput419, keyinput420;
  input keyinput421, keyinput422, keyinput423, keyinput424, keyinput425;
  input keyinput426, keyinput427, keyinput428, keyinput429, keyinput430;
  input keyinput431, keyinput432, keyinput433, keyinput434, keyinput435;

  wire [0:59] keyNTin_Wire_1;
  wire [0:28] KeyNOTWire_1;

  input N26, N189, N138, N68, N143, N91, N159, N101, N219, N156, N116, N72, N90, N121, N246, N135, N86, N42, N130, N13, N195, N29, N106, N75, N87, N8, N85, N126, N51, N259, N152, N55, N171, N73, N165, N177, N201, N153, N1, N74, N80, N261, N237, N146, N96, N268, N59, N17, N89, N88, N111, N149, N36, N255, N267, N228, N207, N210, N183, N260;
  input keyinput256, keyinput257, keyinput258, keyinput259, keyinput260, keyinput261, keyinput262, keyinput263, keyinput264, keyinput265, keyinput266, keyinput267, keyinput268, keyinput269, keyinput270, keyinput271, keyinput272, keyinput273, keyinput274, keyinput275, keyinput276, keyinput277, keyinput278, keyinput279, keyinput280, keyinput281, keyinput282, keyinput283, keyinput284, keyinput285, keyinput286, keyinput287, keyinput288, keyinput289, keyinput290, keyinput291, keyinput292, keyinput293, keyinput294, keyinput295, keyinput296, keyinput297, keyinput298, keyinput299, keyinput300, keyinput301, keyinput302, keyinput303, keyinput304, keyinput305, keyinput306, keyinput307, keyinput308, keyinput309, keyinput310, keyinput311, keyinput312, keyinput313, keyinput314, keyinput315, keyinput316, keyinput317, keyinput318, keyinput319, keyinput320, keyinput321, keyinput322, keyinput323, keyinput324, keyinput325, keyinput326, keyinput327, keyinput328, keyinput329, keyinput330, keyinput331, keyinput332, keyinput333, keyinput334, keyinput335, keyinput336, keyinput337, keyinput338, keyinput339, keyinput340, keyinput341, keyinput342, keyinput343, keyinput344, keyinput345, keyinput346, keyinput347, keyinput348, keyinput349, keyinput350, keyinput351, keyinput352, keyinput353, keyinput354, keyinput355, keyinput356, keyinput357, keyinput358, keyinput359, keyinput360, keyinput361, keyinput362, keyinput363, keyinput364, keyinput365, keyinput366, keyinput367, keyinput368, keyinput369, keyinput370, keyinput371, keyinput372, keyinput373, keyinput374, keyinput375;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83, newWire_84, newWire_85, newWire_86, newWire_87, newWire_88, newWire_89, newWire_90, newWire_91, newWire_92, newWire_93, newWire_94, newWire_95, newWire_96, newWire_97, newWire_98, newWire_99, newWire_100, newWire_101, newWire_102, newWire_103, newWire_104, newWire_105, newWire_106, newWire_107, newWire_108, newWire_109, newWire_110, newWire_111, newWire_112, newWire_113, newWire_114, newWire_115, newWire_116, newWire_117, newWire_118, newWire_119, newWire_120, newWire_121 ;

  xnor KeyGate0 (newWire_0, N26, keyinput256);
  xnor KeyGate1 (newWire_1, N189, keyinput257);
  xor  KeyGate2 (newWire_2, N138, keyinput258);
  xor  KeyGate3 (keyNTin_Wire_1[0], N68, keyinput259);
  xnor keyNTinGate_1_0(KeyNOTWire_1[0], keyinput376, keyNTin_Wire_1[0]);
  not KeyNOTGate_1_0(newWire_3, KeyNOTWire_1[0]);
  xor  KeyGate4 (keyNTin_Wire_1[1], N143, keyinput260);
  xor keyNTinGate_1_1(KeyNOTWire_1[1], keyinput377, keyNTin_Wire_1[1]);
  not KeyNOTGate_1_1(newWire_4, KeyNOTWire_1[1]);
  xor  KeyGate5 (keyNTin_Wire_1[2], N91, keyinput261);
  xnor keyNTinGate_1_2(KeyNOTWire_1[2], keyinput378, keyNTin_Wire_1[2]);
  not KeyNOTGate_1_2(newWire_5, KeyNOTWire_1[2]);
  xor  KeyGate6 (newWire_6, N159, keyinput262);
  xor  KeyGate7 (newWire_7, N101, keyinput263);
  xor  KeyGate8 (newWire_8, N219, keyinput264);
  xnor KeyGate9 (newWire_9, N156, keyinput265);
  xnor KeyGate10 (keyNTin_Wire_1[3], N116, keyinput266);
  xor keyNTinGate_1_3(newWire_10, keyinput379, keyNTin_Wire_1[3]);
  xor  KeyGate11 (keyNTin_Wire_1[4], N72, keyinput267);
  xnor keyNTinGate_1_4(KeyNOTWire_1[3], keyinput380, keyNTin_Wire_1[4]);
  not KeyNOTGate_1_3(newWire_11, KeyNOTWire_1[3]);
  xnor KeyGate12 (newWire_12, N90, keyinput268);
  xnor KeyGate13 (keyNTin_Wire_1[5], N121, keyinput269);
  xnor keyNTinGate_1_5(newWire_13, keyinput381, keyNTin_Wire_1[5]);
  xnor KeyGate14 (keyNTin_Wire_1[6], N246, keyinput270);
  xnor keyNTinGate_1_6(KeyNOTWire_1[4], keyinput382, keyNTin_Wire_1[6]);
  not KeyNOTGate_1_4(newWire_14, KeyNOTWire_1[4]);
  xor  KeyGate15 (keyNTin_Wire_1[7], N135, keyinput271);
  xor keyNTinGate_1_7(KeyNOTWire_1[5], keyinput383, keyNTin_Wire_1[7]);
  not KeyNOTGate_1_5(newWire_15, KeyNOTWire_1[5]);
  xor  KeyGate16 (keyNTin_Wire_1[8], N86, keyinput272);
  xnor keyNTinGate_1_8(KeyNOTWire_1[6], keyinput384, keyNTin_Wire_1[8]);
  not KeyNOTGate_1_6(newWire_16, KeyNOTWire_1[6]);
  xnor KeyGate17 (keyNTin_Wire_1[9], N42, keyinput273);
  xor keyNTinGate_1_9(newWire_17, keyinput385, keyNTin_Wire_1[9]);
  xnor KeyGate18 (newWire_18, N130, keyinput274);
  xor  KeyGate19 (newWire_19, N13, keyinput275);
  xor  KeyGate20 (newWire_20, N195, keyinput276);
  xor  KeyGate21 (newWire_21, N29, keyinput277);
  xnor KeyGate22 (newWire_22, N106, keyinput278);
  xnor KeyGate23 (keyNTin_Wire_1[10], N75, keyinput279);
  xnor keyNTinGate_1_10(KeyNOTWire_1[7], keyinput386, keyNTin_Wire_1[10]);
  not KeyNOTGate_1_7(newWire_23, KeyNOTWire_1[7]);
  xor  KeyGate24 (newWire_24, N87, keyinput280);
  xor  KeyGate25 (keyNTin_Wire_1[11], N8, keyinput281);
  xor keyNTinGate_1_11(newWire_25, keyinput387, keyNTin_Wire_1[11]);
  xnor KeyGate26 (newWire_26, N85, keyinput282);
  xnor KeyGate27 (keyNTin_Wire_1[12], N126, keyinput283);
  xor keyNTinGate_1_12(newWire_27, keyinput388, keyNTin_Wire_1[12]);
  xnor KeyGate28 (newWire_28, N51, keyinput284);
  xnor KeyGate29 (newWire_29, N259, keyinput285);
  xnor KeyGate30 (newWire_30, N152, keyinput286);
  xnor KeyGate31 (newWire_31, N55, keyinput287);
  xnor KeyGate32 (keyNTin_Wire_1[13], N171, keyinput288);
  xnor keyNTinGate_1_13(KeyNOTWire_1[8], keyinput389, keyNTin_Wire_1[13]);
  not KeyNOTGate_1_8(newWire_32, KeyNOTWire_1[8]);
  xor  KeyGate33 (newWire_33, N73, keyinput289);
  xor  KeyGate34 (keyNTin_Wire_1[14], N165, keyinput290);
  xor keyNTinGate_1_14(KeyNOTWire_1[9], keyinput390, keyNTin_Wire_1[14]);
  not KeyNOTGate_1_9(newWire_34, KeyNOTWire_1[9]);
  xor  KeyGate35 (keyNTin_Wire_1[15], N177, keyinput291);
  xor keyNTinGate_1_15(newWire_35, keyinput391, keyNTin_Wire_1[15]);
  xor  KeyGate36 (keyNTin_Wire_1[16], N201, keyinput292);
  xnor keyNTinGate_1_16(newWire_36, keyinput392, keyNTin_Wire_1[16]);
  xor  KeyGate37 (keyNTin_Wire_1[17], N153, keyinput293);
  xor keyNTinGate_1_17(newWire_37, keyinput393, keyNTin_Wire_1[17]);
  xnor KeyGate38 (newWire_38, N1, keyinput294);
  xnor KeyGate39 (newWire_39, N74, keyinput295);
  xnor KeyGate40 (keyNTin_Wire_1[18], N80, keyinput296);
  xnor keyNTinGate_1_18(newWire_40, keyinput394, keyNTin_Wire_1[18]);
  xor  KeyGate41 (keyNTin_Wire_1[19], N261, keyinput297);
  xnor keyNTinGate_1_19(KeyNOTWire_1[10], keyinput395, keyNTin_Wire_1[19]);
  not KeyNOTGate_1_10(newWire_41, KeyNOTWire_1[10]);
  xnor KeyGate42 (keyNTin_Wire_1[20], N237, keyinput298);
  xor keyNTinGate_1_20(KeyNOTWire_1[11], keyinput396, keyNTin_Wire_1[20]);
  not KeyNOTGate_1_11(newWire_42, KeyNOTWire_1[11]);
  xnor KeyGate43 (newWire_43, N146, keyinput299);
  xnor KeyGate44 (newWire_44, N96, keyinput300);
  xor  KeyGate45 (keyNTin_Wire_1[21], N268, keyinput301);
  xor keyNTinGate_1_21(newWire_45, keyinput397, keyNTin_Wire_1[21]);
  xnor KeyGate46 (keyNTin_Wire_1[22], N59, keyinput302);
  xnor keyNTinGate_1_22(KeyNOTWire_1[12], keyinput398, keyNTin_Wire_1[22]);
  not KeyNOTGate_1_12(newWire_46, KeyNOTWire_1[12]);
  xor  KeyGate47 (keyNTin_Wire_1[23], N17, keyinput303);
  xor keyNTinGate_1_23(KeyNOTWire_1[13], keyinput399, keyNTin_Wire_1[23]);
  not KeyNOTGate_1_13(newWire_47, KeyNOTWire_1[13]);
  xor  KeyGate48 (keyNTin_Wire_1[24], N89, keyinput304);
  xnor keyNTinGate_1_24(KeyNOTWire_1[14], keyinput400, keyNTin_Wire_1[24]);
  not KeyNOTGate_1_14(newWire_48, KeyNOTWire_1[14]);
  xor  KeyGate49 (keyNTin_Wire_1[25], N88, keyinput305);
  xor keyNTinGate_1_25(newWire_49, keyinput401, keyNTin_Wire_1[25]);
  xor  KeyGate50 (keyNTin_Wire_1[26], N111, keyinput306);
  xnor keyNTinGate_1_26(newWire_50, keyinput402, keyNTin_Wire_1[26]);
  xor  KeyGate51 (keyNTin_Wire_1[27], N149, keyinput307);
  xnor keyNTinGate_1_27(KeyNOTWire_1[15], keyinput403, keyNTin_Wire_1[27]);
  not KeyNOTGate_1_15(newWire_51, KeyNOTWire_1[15]);
  xor  KeyGate52 (newWire_52, N36, keyinput308);
  xnor KeyGate53 (keyNTin_Wire_1[28], N255, keyinput309);
  xor keyNTinGate_1_28(KeyNOTWire_1[16], keyinput404, keyNTin_Wire_1[28]);
  not KeyNOTGate_1_16(newWire_53, KeyNOTWire_1[16]);
  xor  KeyGate54 (keyNTin_Wire_1[29], N267, keyinput310);
  xnor keyNTinGate_1_29(newWire_54, keyinput405, keyNTin_Wire_1[29]);
  xnor KeyGate55 (newWire_55, N228, keyinput311);
  xnor KeyGate56 (newWire_56, N207, keyinput312);
  xnor KeyGate57 (newWire_57, N210, keyinput313);
  xnor KeyGate58 (newWire_58, N183, keyinput314);
  xor  KeyGate59 (keyNTin_Wire_1[30], N260, keyinput315);
  xnor keyNTinGate_1_30(KeyNOTWire_1[17], keyinput406, keyNTin_Wire_1[30]);
  not KeyNOTGate_1_17(newWire_59, KeyNOTWire_1[17]);
  xor  KeyGate60 (newWire_60, N26, keyinput316);
  xnor KeyGate61 (newWire_61, N189, keyinput317);
  xor  KeyGate62 (keyNTin_Wire_1[31], N138, keyinput318);
  xnor keyNTinGate_1_31(newWire_62, keyinput407, keyNTin_Wire_1[31]);
  xnor KeyGate63 (newWire_63, N68, keyinput319);
  xnor KeyGate64 (newWire_64, N143, keyinput320);
  xnor KeyGate65 (keyNTin_Wire_1[32], N91, keyinput321);
  xnor keyNTinGate_1_32(newWire_65, keyinput408, keyNTin_Wire_1[32]);
  xor  KeyGate66 (keyNTin_Wire_1[33], N159, keyinput322);
  xor keyNTinGate_1_33(newWire_66, keyinput409, keyNTin_Wire_1[33]);
  xor  KeyGate67 (newWire_67, N101, keyinput323);
  xor  KeyGate68 (keyNTin_Wire_1[34], N219, keyinput324);
  xor keyNTinGate_1_34(KeyNOTWire_1[18], keyinput410, keyNTin_Wire_1[34]);
  not KeyNOTGate_1_18(newWire_68, KeyNOTWire_1[18]);
  xor  KeyGate69 (newWire_69, N156, keyinput325);
  xnor KeyGate70 (keyNTin_Wire_1[35], N116, keyinput326);
  xnor keyNTinGate_1_35(KeyNOTWire_1[19], keyinput411, keyNTin_Wire_1[35]);
  not KeyNOTGate_1_19(newWire_70, KeyNOTWire_1[19]);
  xor  KeyGate71 (newWire_71, N72, keyinput327);
  xor  KeyGate72 (newWire_72, N90, keyinput328);
  xor  KeyGate73 (newWire_73, N121, keyinput329);
  xnor KeyGate74 (keyNTin_Wire_1[36], N246, keyinput330);
  xor keyNTinGate_1_36(KeyNOTWire_1[20], keyinput412, keyNTin_Wire_1[36]);
  not KeyNOTGate_1_20(newWire_74, KeyNOTWire_1[20]);
  xnor KeyGate75 (keyNTin_Wire_1[37], N135, keyinput331);
  xor keyNTinGate_1_37(KeyNOTWire_1[21], keyinput413, keyNTin_Wire_1[37]);
  not KeyNOTGate_1_21(newWire_75, KeyNOTWire_1[21]);
  xnor KeyGate76 (newWire_76, N86, keyinput332);
  xnor KeyGate77 (keyNTin_Wire_1[38], N42, keyinput333);
  xor keyNTinGate_1_38(newWire_77, keyinput414, keyNTin_Wire_1[38]);
  xor  KeyGate78 (newWire_78, N130, keyinput334);
  xnor KeyGate79 (newWire_79, N13, keyinput335);
  xnor KeyGate80 (newWire_80, N195, keyinput336);
  xnor KeyGate81 (keyNTin_Wire_1[39], N29, keyinput337);
  xor keyNTinGate_1_39(newWire_81, keyinput415, keyNTin_Wire_1[39]);
  xnor KeyGate82 (newWire_82, N106, keyinput338);
  xnor KeyGate83 (keyNTin_Wire_1[40], N75, keyinput339);
  xor keyNTinGate_1_40(KeyNOTWire_1[22], keyinput416, keyNTin_Wire_1[40]);
  not KeyNOTGate_1_22(newWire_83, KeyNOTWire_1[22]);
  xnor KeyGate84 (newWire_84, N87, keyinput340);
  xor  KeyGate85 (keyNTin_Wire_1[41], N8, keyinput341);
  xor keyNTinGate_1_41(KeyNOTWire_1[23], keyinput417, keyNTin_Wire_1[41]);
  not KeyNOTGate_1_23(newWire_85, KeyNOTWire_1[23]);
  xnor KeyGate86 (newWire_86, N85, keyinput342);
  xnor KeyGate87 (newWire_87, N126, keyinput343);
  xnor KeyGate88 (newWire_88, N51, keyinput344);
  xnor KeyGate89 (newWire_89, N259, keyinput345);
  xnor KeyGate90 (keyNTin_Wire_1[42], N152, keyinput346);
  xnor keyNTinGate_1_42(KeyNOTWire_1[24], keyinput418, keyNTin_Wire_1[42]);
  not KeyNOTGate_1_24(newWire_90, KeyNOTWire_1[24]);
  xnor KeyGate91 (keyNTin_Wire_1[43], N55, keyinput347);
  xnor keyNTinGate_1_43(newWire_91, keyinput419, keyNTin_Wire_1[43]);
  xor  KeyGate92 (newWire_92, N171, keyinput348);
  xor  KeyGate93 (keyNTin_Wire_1[44], N73, keyinput349);
  xor keyNTinGate_1_44(newWire_93, keyinput420, keyNTin_Wire_1[44]);
  xnor KeyGate94 (newWire_94, N165, keyinput350);
  xor  KeyGate95 (newWire_95, N177, keyinput351);
  xnor KeyGate96 (keyNTin_Wire_1[45], N201, keyinput352);
  xor keyNTinGate_1_45(newWire_96, keyinput421, keyNTin_Wire_1[45]);
  xor  KeyGate97 (keyNTin_Wire_1[46], N153, keyinput353);
  xor keyNTinGate_1_46(newWire_97, keyinput422, keyNTin_Wire_1[46]);
  xor  KeyGate98 (keyNTin_Wire_1[47], N1, keyinput354);
  xnor keyNTinGate_1_47(KeyNOTWire_1[25], keyinput423, keyNTin_Wire_1[47]);
  not KeyNOTGate_1_25(newWire_98, KeyNOTWire_1[25]);
  xnor KeyGate99 (keyNTin_Wire_1[48], N74, keyinput355);
  xnor keyNTinGate_1_48(newWire_99, keyinput424, keyNTin_Wire_1[48]);
  xor  KeyGate100 (newWire_100, N80, keyinput356);
  xor  KeyGate101 (newWire_101, N261, keyinput357);
  xor  KeyGate102 (keyNTin_Wire_1[49], N237, keyinput358);
  xnor keyNTinGate_1_49(newWire_102, keyinput425, keyNTin_Wire_1[49]);
  xor  KeyGate103 (newWire_103, N146, keyinput359);
  xnor KeyGate104 (newWire_104, N96, keyinput360);
  xnor KeyGate105 (newWire_105, N268, keyinput361);
  xnor KeyGate106 (keyNTin_Wire_1[50], N59, keyinput362);
  xor keyNTinGate_1_50(newWire_106, keyinput426, keyNTin_Wire_1[50]);
  xor  KeyGate107 (keyNTin_Wire_1[51], N17, keyinput363);
  xnor keyNTinGate_1_51(KeyNOTWire_1[26], keyinput427, keyNTin_Wire_1[51]);
  not KeyNOTGate_1_26(newWire_107, KeyNOTWire_1[26]);
  xor  KeyGate108 (keyNTin_Wire_1[52], N89, keyinput364);
  xnor keyNTinGate_1_52(KeyNOTWire_1[27], keyinput428, keyNTin_Wire_1[52]);
  not KeyNOTGate_1_27(newWire_108, KeyNOTWire_1[27]);
  xor  KeyGate109 (keyNTin_Wire_1[53], N88, keyinput365);
  xnor keyNTinGate_1_53(newWire_109, keyinput429, keyNTin_Wire_1[53]);
  xor  KeyGate110 (newWire_110, N111, keyinput366);
  xnor KeyGate111 (newWire_111, N149, keyinput367);
  xnor KeyGate112 (keyNTin_Wire_1[54], N36, keyinput368);
  xor keyNTinGate_1_54(newWire_112, keyinput430, keyNTin_Wire_1[54]);
  xor  KeyGate113 (keyNTin_Wire_1[55], N255, keyinput369);
  xor keyNTinGate_1_55(KeyNOTWire_1[28], keyinput431, keyNTin_Wire_1[55]);
  not KeyNOTGate_1_28(newWire_113, KeyNOTWire_1[28]);
  xor  KeyGate114 (newWire_114, N267, keyinput370);
  xnor KeyGate115 (newWire_115, N228, keyinput371);
  xnor KeyGate116 (newWire_116, N207, keyinput372);
  xnor KeyGate117 (keyNTin_Wire_1[56], N210, keyinput373);
  xnor keyNTinGate_1_56(newWire_117, keyinput432, keyNTin_Wire_1[56]);
  xor  KeyGate118 (newWire_118, N183, keyinput374);
  xnor KeyGate119 (newWire_119, N260, keyinput375);
  and some_function (keyNTin_Wire_1[57], newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59 );
  xor keyNTinGate_1_57(newWire_120, keyinput433, keyNTin_Wire_1[57]);
  nand compl_function (keyNTin_Wire_1[58], newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83, newWire_84, newWire_85, newWire_86, newWire_87, newWire_88, newWire_89, newWire_90, newWire_91, newWire_92, newWire_93, newWire_94, newWire_95, newWire_96, newWire_97, newWire_98, newWire_99, newWire_100, newWire_101, newWire_102, newWire_103, newWire_104, newWire_105, newWire_106, newWire_107, newWire_108, newWire_109, newWire_110, newWire_111, newWire_112, newWire_113, newWire_114, newWire_115, newWire_116, newWire_117, newWire_118, newWire_119);
  xor keyNTinGate_1_58(newWire_121, keyinput434, keyNTin_Wire_1[58]);
  and finalAND (keyNTin_Wire_1[59], newWire_120, newWire_121);
  xnor keyNTinGate_1_59(KeyWire_0_2, keyinput435, keyNTin_Wire_1[59]);

endmodule /* AntiSAT */
