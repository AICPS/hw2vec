`timescale 1ns / 1ps
// Verilog
// c499
// Ninputs 41
// Noutputs 32
// NtotalGates 202
// XOR2 104
// AND2 40
// NOT1 40
// AND4 8
// OR4 2
// AND5 8

module top (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
                  N753,N754,N755,
        keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4,
        keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9,
        keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14,
        keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19,
        keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24,
        keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29,
        keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34,
        keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39,
        keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44,
        keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49,
        keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54,
        keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59,
        keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63);

  input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4;
  input keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9;
  input keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14;
  input keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19;
  input keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24;
  input keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29;
  input keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34;
  input keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39;
  input keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44;
  input keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49;
  input keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54;
  input keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59;
  input keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63;

  wire [0:63] KeyWire_0;
  wire [0:34] KeyNOTWire_0;

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;

output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723;

xor XOR2_1 (N250, N1, N5);
xor XOR2_2 (N251, N9, N13);
xor XOR2_3 (N252, N17, N21);
  xor XOR2_4 (KeyWire_0[0], N25, N29);
  xnor KeyGate_0_0(KeyNOTWire_0[0], keyIn_0_0, KeyWire_0[0]);
  not KeyNOTGate_0_0(N253, KeyNOTWire_0[0]);
  xor XOR2_5 (KeyWire_0[1], N33, N37);
  xnor KeyGate_0_1(KeyNOTWire_0[1], keyIn_0_1, KeyWire_0[1]);
  not KeyNOTGate_0_1(N254, KeyNOTWire_0[1]);
  xor XOR2_6 (KeyWire_0[2], N41, N45);
  xor KeyGate_0_2(N255, keyIn_0_2, KeyWire_0[2]);
  xor XOR2_7 (KeyWire_0[3], N49, N53);
  xnor KeyGate_0_3(N256, keyIn_0_3, KeyWire_0[3]);
  xor XOR2_8 (KeyWire_0[4], N57, N61);
  xnor KeyGate_0_4(N257, keyIn_0_4, KeyWire_0[4]);
  xor XOR2_9 (KeyWire_0[5], N65, N69);
  xor KeyGate_0_5(N258, keyIn_0_5, KeyWire_0[5]);
xor XOR2_10 (N259, N73, N77);
xor XOR2_11 (N260, N81, N85);
xor XOR2_12 (N261, N89, N93);
xor XOR2_13 (N262, N97, N101);
xor XOR2_14 (N263, N105, N109);
xor XOR2_15 (N264, N113, N117);
xor XOR2_16 (N265, N121, N125);
and AND2_17 (N266, N129, N137);
and AND2_18 (N267, N130, N137);
and AND2_19 (N268, N131, N137);
and AND2_20 (N269, N132, N137);
and AND2_21 (N270, N133, N137);
and AND2_22 (N271, N134, N137);
and AND2_23 (N272, N135, N137);
and AND2_24 (N273, N136, N137);
xor XOR2_25 (N274, N1, N17);
xor XOR2_26 (N275, N33, N49);
xor XOR2_27 (N276, N5, N21);
xor XOR2_28 (N277, N37, N53);
xor XOR2_29 (N278, N9, N25);
xor XOR2_30 (N279, N41, N57);
xor XOR2_31 (N280, N13, N29);
xor XOR2_32 (N281, N45, N61);
xor XOR2_33 (N282, N65, N81);
xor XOR2_34 (N283, N97, N113);
xor XOR2_35 (N284, N69, N85);
xor XOR2_36 (N285, N101, N117);
xor XOR2_37 (N286, N73, N89);
xor XOR2_38 (N287, N105, N121);
xor XOR2_39 (N288, N77, N93);
xor XOR2_40 (N289, N109, N125);
  xor XOR2_41 (KeyWire_0[6], N250, N251);
  xnor KeyGate_0_6(KeyNOTWire_0[2], keyIn_0_6, KeyWire_0[6]);
  not KeyNOTGate_0_2(N290, KeyNOTWire_0[2]);
  xor XOR2_42 (KeyWire_0[7], N252, N253);
  xnor KeyGate_0_7(N293, keyIn_0_7, KeyWire_0[7]);
  xor XOR2_43 (KeyWire_0[8], N254, N255);
  xor KeyGate_0_8(KeyNOTWire_0[3], keyIn_0_8, KeyWire_0[8]);
  not KeyNOTGate_0_3(N296, KeyNOTWire_0[3]);
  xor XOR2_44 (KeyWire_0[9], N256, N257);
  xnor KeyGate_0_9(N299, keyIn_0_9, KeyWire_0[9]);
  xor XOR2_45 (KeyWire_0[10], N258, N259);
  xnor KeyGate_0_10(N302, keyIn_0_10, KeyWire_0[10]);
  xor XOR2_46 (KeyWire_0[11], N260, N261);
  xnor KeyGate_0_11(KeyNOTWire_0[4], keyIn_0_11, KeyWire_0[11]);
  not KeyNOTGate_0_4(N305, KeyNOTWire_0[4]);
  xor XOR2_47 (KeyWire_0[12], N262, N263);
  xor KeyGate_0_12(KeyNOTWire_0[5], keyIn_0_12, KeyWire_0[12]);
  not KeyNOTGate_0_5(N308, KeyNOTWire_0[5]);
  xor XOR2_48 (KeyWire_0[13], N264, N265);
  xor KeyGate_0_13(KeyNOTWire_0[6], keyIn_0_13, KeyWire_0[13]);
  not KeyNOTGate_0_6(N311, KeyNOTWire_0[6]);
  xor XOR2_49 (KeyWire_0[14], N274, N275);
  xor KeyGate_0_14(KeyNOTWire_0[7], keyIn_0_14, KeyWire_0[14]);
  not KeyNOTGate_0_7(N314, KeyNOTWire_0[7]);
  xor XOR2_50 (KeyWire_0[15], N276, N277);
  xnor KeyGate_0_15(KeyNOTWire_0[8], keyIn_0_15, KeyWire_0[15]);
  not KeyNOTGate_0_8(N315, KeyNOTWire_0[8]);
  xor XOR2_51 (KeyWire_0[16], N278, N279);
  xnor KeyGate_0_16(KeyNOTWire_0[9], keyIn_0_16, KeyWire_0[16]);
  not KeyNOTGate_0_9(N316, KeyNOTWire_0[9]);
  xor XOR2_52 (KeyWire_0[17], N280, N281);
  xor KeyGate_0_17(N317, keyIn_0_17, KeyWire_0[17]);
  xor XOR2_53 (KeyWire_0[18], N282, N283);
  xor KeyGate_0_18(N318, keyIn_0_18, KeyWire_0[18]);
  xor XOR2_54 (KeyWire_0[19], N284, N285);
  xnor KeyGate_0_19(N319, keyIn_0_19, KeyWire_0[19]);
  xor XOR2_55 (KeyWire_0[20], N286, N287);
  xor KeyGate_0_20(KeyNOTWire_0[10], keyIn_0_20, KeyWire_0[20]);
  not KeyNOTGate_0_10(N320, KeyNOTWire_0[10]);
  xor XOR2_56 (KeyWire_0[21], N288, N289);
  xnor KeyGate_0_21(KeyNOTWire_0[11], keyIn_0_21, KeyWire_0[21]);
  not KeyNOTGate_0_11(N321, KeyNOTWire_0[11]);
  xor XOR2_57 (KeyWire_0[22], N290, N293);
  xnor KeyGate_0_22(KeyNOTWire_0[12], keyIn_0_22, KeyWire_0[22]);
  not KeyNOTGate_0_12(N338, KeyNOTWire_0[12]);
  xor XOR2_58 (KeyWire_0[23], N296, N299);
  xnor KeyGate_0_23(N339, keyIn_0_23, KeyWire_0[23]);
  xor XOR2_59 (KeyWire_0[24], N290, N296);
  xor KeyGate_0_24(KeyNOTWire_0[13], keyIn_0_24, KeyWire_0[24]);
  not KeyNOTGate_0_13(N340, KeyNOTWire_0[13]);
  xor XOR2_60 (KeyWire_0[25], N293, N299);
  xor KeyGate_0_25(KeyNOTWire_0[14], keyIn_0_25, KeyWire_0[25]);
  not KeyNOTGate_0_14(N341, KeyNOTWire_0[14]);
  xor XOR2_61 (KeyWire_0[26], N302, N305);
  xor KeyGate_0_26(N342, keyIn_0_26, KeyWire_0[26]);
  xor XOR2_62 (KeyWire_0[27], N308, N311);
  xor KeyGate_0_27(N343, keyIn_0_27, KeyWire_0[27]);
  xor XOR2_63 (KeyWire_0[28], N302, N308);
  xnor KeyGate_0_28(N344, keyIn_0_28, KeyWire_0[28]);
  xor XOR2_64 (KeyWire_0[29], N305, N311);
  xnor KeyGate_0_29(N345, keyIn_0_29, KeyWire_0[29]);
  xor XOR2_65 (KeyWire_0[30], N266, N342);
  xor KeyGate_0_30(KeyNOTWire_0[15], keyIn_0_30, KeyWire_0[30]);
  not KeyNOTGate_0_15(N346, KeyNOTWire_0[15]);
  xor XOR2_66 (KeyWire_0[31], N267, N343);
  xor KeyGate_0_31(KeyNOTWire_0[16], keyIn_0_31, KeyWire_0[31]);
  not KeyNOTGate_0_16(N347, KeyNOTWire_0[16]);
  xor XOR2_67 (KeyWire_0[32], N268, N344);
  xor KeyGate_0_32(KeyNOTWire_0[17], keyIn_0_32, KeyWire_0[32]);
  not KeyNOTGate_0_17(N348, KeyNOTWire_0[17]);
  xor XOR2_68 (KeyWire_0[33], N269, N345);
  xor KeyGate_0_33(N349, keyIn_0_33, KeyWire_0[33]);
  xor XOR2_69 (KeyWire_0[34], N270, N338);
  xnor KeyGate_0_34(KeyNOTWire_0[18], keyIn_0_34, KeyWire_0[34]);
  not KeyNOTGate_0_18(N350, KeyNOTWire_0[18]);
  xor XOR2_70 (KeyWire_0[35], N271, N339);
  xor KeyGate_0_35(N351, keyIn_0_35, KeyWire_0[35]);
  xor XOR2_71 (KeyWire_0[36], N272, N340);
  xnor KeyGate_0_36(KeyNOTWire_0[19], keyIn_0_36, KeyWire_0[36]);
  not KeyNOTGate_0_19(N352, KeyNOTWire_0[19]);
  xor XOR2_72 (KeyWire_0[37], N273, N341);
  xor KeyGate_0_37(N353, keyIn_0_37, KeyWire_0[37]);
  xor XOR2_73 (KeyWire_0[38], N314, N346);
  xnor KeyGate_0_38(N354, keyIn_0_38, KeyWire_0[38]);
  xor XOR2_74 (KeyWire_0[39], N315, N347);
  xor KeyGate_0_39(KeyNOTWire_0[20], keyIn_0_39, KeyWire_0[39]);
  not KeyNOTGate_0_20(N367, KeyNOTWire_0[20]);
  xor XOR2_75 (KeyWire_0[40], N316, N348);
  xnor KeyGate_0_40(KeyNOTWire_0[21], keyIn_0_40, KeyWire_0[40]);
  not KeyNOTGate_0_21(N380, KeyNOTWire_0[21]);
  xor XOR2_76 (KeyWire_0[41], N317, N349);
  xor KeyGate_0_41(KeyNOTWire_0[22], keyIn_0_41, KeyWire_0[41]);
  not KeyNOTGate_0_22(N393, KeyNOTWire_0[22]);
  xor XOR2_77 (KeyWire_0[42], N318, N350);
  xnor KeyGate_0_42(N406, keyIn_0_42, KeyWire_0[42]);
  xor XOR2_78 (KeyWire_0[43], N319, N351);
  xnor KeyGate_0_43(N419, keyIn_0_43, KeyWire_0[43]);
  xor XOR2_79 (KeyWire_0[44], N320, N352);
  xor KeyGate_0_44(KeyNOTWire_0[23], keyIn_0_44, KeyWire_0[44]);
  not KeyNOTGate_0_23(N432, KeyNOTWire_0[23]);
  xor XOR2_80 (KeyWire_0[45], N321, N353);
  xnor KeyGate_0_45(KeyNOTWire_0[24], keyIn_0_45, KeyWire_0[45]);
  not KeyNOTGate_0_24(N445, KeyNOTWire_0[24]);
not NOT1_81 (N554, N354);
not NOT1_82 (N555, N367);
not NOT1_83 (N556, N380);
not NOT1_84 (N557, N354);
not NOT1_85 (N558, N367);
not NOT1_86 (N559, N393);
not NOT1_87 (N560, N354);
not NOT1_88 (N561, N380);
not NOT1_89 (N562, N393);
not NOT1_90 (N563, N367);
not NOT1_91 (N564, N380);
not NOT1_92 (N565, N393);
not NOT1_93 (N566, N419);
not NOT1_94 (N567, N445);
not NOT1_95 (N568, N419);
not NOT1_96 (N569, N432);
not NOT1_97 (N570, N406);
not NOT1_98 (N571, N445);
not NOT1_99 (N572, N406);
not NOT1_100 (N573, N432);
not NOT1_101 (N574, N406);
not NOT1_102 (N575, N419);
not NOT1_103 (N576, N432);
not NOT1_104 (N577, N406);
not NOT1_105 (N578, N419);
not NOT1_106 (N579, N445);
not NOT1_107 (N580, N406);
not NOT1_108 (N581, N432);
not NOT1_109 (N582, N445);
not NOT1_110 (N583, N419);
not NOT1_111 (N584, N432);
not NOT1_112 (N585, N445);
not NOT1_113 (N586, N367);
not NOT1_114 (N587, N393);
not NOT1_115 (N588, N367);
not NOT1_116 (N589, N380);
not NOT1_117 (N590, N354);
not NOT1_118 (N591, N393);
not NOT1_119 (N592, N354);
not NOT1_120 (N593, N380);
  and AND4_121 (KeyWire_0[46], N554, N555, N556, N393);
  xor KeyGate_0_46(KeyNOTWire_0[25], keyIn_0_46, KeyWire_0[46]);
  not KeyNOTGate_0_25(N594, KeyNOTWire_0[25]);
  and AND4_122 (KeyWire_0[47], N557, N558, N380, N559);
  xnor KeyGate_0_47(KeyNOTWire_0[26], keyIn_0_47, KeyWire_0[47]);
  not KeyNOTGate_0_26(N595, KeyNOTWire_0[26]);
  and AND4_123 (KeyWire_0[48], N560, N367, N561, N562);
  xnor KeyGate_0_48(N596, keyIn_0_48, KeyWire_0[48]);
  and AND4_124 (KeyWire_0[49], N354, N563, N564, N565);
  xnor KeyGate_0_49(KeyNOTWire_0[27], keyIn_0_49, KeyWire_0[49]);
  not KeyNOTGate_0_27(N597, KeyNOTWire_0[27]);
  and AND4_125 (KeyWire_0[50], N574, N575, N576, N445);
  xnor KeyGate_0_50(KeyNOTWire_0[28], keyIn_0_50, KeyWire_0[50]);
  not KeyNOTGate_0_28(N598, KeyNOTWire_0[28]);
  and AND4_126 (KeyWire_0[51], N577, N578, N432, N579);
  xnor KeyGate_0_51(N599, keyIn_0_51, KeyWire_0[51]);
  and AND4_127 (KeyWire_0[52], N580, N419, N581, N582);
  xnor KeyGate_0_52(KeyNOTWire_0[29], keyIn_0_52, KeyWire_0[52]);
  not KeyNOTGate_0_29(N600, KeyNOTWire_0[29]);
  and AND4_128 (KeyWire_0[53], N406, N583, N584, N585);
  xor KeyGate_0_53(KeyNOTWire_0[30], keyIn_0_53, KeyWire_0[53]);
  not KeyNOTGate_0_30(N601, KeyNOTWire_0[30]);
  or OR4_129 (KeyWire_0[54], N594, N595, N596, N597);
  xnor KeyGate_0_54(KeyNOTWire_0[31], keyIn_0_54, KeyWire_0[54]);
  not KeyNOTGate_0_31(N602, KeyNOTWire_0[31]);
  or OR4_130 (KeyWire_0[55], N598, N599, N600, N601);
  xor KeyGate_0_55(N607, keyIn_0_55, KeyWire_0[55]);
  and AND5_131 (KeyWire_0[56], N406, N566, N432, N567, N602);
  xnor KeyGate_0_56(N620, keyIn_0_56, KeyWire_0[56]);
  and AND5_132 (KeyWire_0[57], N406, N568, N569, N445, N602);
  xnor KeyGate_0_57(N625, keyIn_0_57, KeyWire_0[57]);
  and AND5_133 (KeyWire_0[58], N570, N419, N432, N571, N602);
  xor KeyGate_0_58(KeyNOTWire_0[32], keyIn_0_58, KeyWire_0[58]);
  not KeyNOTGate_0_32(N630, KeyNOTWire_0[32]);
  and AND5_134 (KeyWire_0[59], N572, N419, N573, N445, N602);
  xnor KeyGate_0_59(N635, keyIn_0_59, KeyWire_0[59]);
  and AND5_135 (KeyWire_0[60], N354, N586, N380, N587, N607);
  xnor KeyGate_0_60(KeyNOTWire_0[33], keyIn_0_60, KeyWire_0[60]);
  not KeyNOTGate_0_33(N640, KeyNOTWire_0[33]);
  and AND5_136 (KeyWire_0[61], N354, N588, N589, N393, N607);
  xor KeyGate_0_61(N645, keyIn_0_61, KeyWire_0[61]);
  and AND5_137 (KeyWire_0[62], N590, N367, N380, N591, N607);
  xnor KeyGate_0_62(KeyNOTWire_0[34], keyIn_0_62, KeyWire_0[62]);
  not KeyNOTGate_0_34(N650, KeyNOTWire_0[34]);
  and AND5_138 (KeyWire_0[63], N592, N367, N593, N393, N607);
  xor KeyGate_0_63(N655, keyIn_0_63, KeyWire_0[63]);
and AND2_139 (N692, N354, N620);
and AND2_140 (N693, N367, N620);
and AND2_141 (N694, N380, N620);
and AND2_142 (N695, N393, N620);
and AND2_143 (N696, N354, N625);
and AND2_144 (N697, N367, N625);
and AND2_145 (N698, N380, N625);
and AND2_146 (N699, N393, N625);
and AND2_147 (N700, N354, N630);
and AND2_148 (N701, N367, N630);
and AND2_149 (N702, N380, N630);
and AND2_150 (N703, N393, N630);
and AND2_151 (N704, N354, N635);
and AND2_152 (N705, N367, N635);
and AND2_153 (N706, N380, N635);
and AND2_154 (N707, N393, N635);
and AND2_155 (N708, N406, N640);
and AND2_156 (N709, N419, N640);
and AND2_157 (N710, N432, N640);
and AND2_158 (N711, N445, N640);
and AND2_159 (N712, N406, N645);
and AND2_160 (N713, N419, N645);
and AND2_161 (N714, N432, N645);
and AND2_162 (N715, N445, N645);
and AND2_163 (N716, N406, N650);
and AND2_164 (N717, N419, N650);
and AND2_165 (N718, N432, N650);
and AND2_166 (N719, N445, N650);
and AND2_167 (N720, N406, N655);
and AND2_168 (N721, N419, N655);
and AND2_169 (N722, N432, N655);
and AND2_170 (N723, N445, N655);
xor XOR2_171 (N724, N1, N692);
xor XOR2_172 (N725, N5, N693);
xor XOR2_173 (N726, N9, N694);
xor XOR2_174 (N727, N13, N695);
xor XOR2_175 (N728, N17, N696);
xor XOR2_176 (N729, N21, N697);
xor XOR2_177 (N730, N25, N698);
xor XOR2_178 (N731, N29, N699);
xor XOR2_179 (N732, N33, N700);
xor XOR2_180 (N733, N37, N701);
xor XOR2_181 (N734, N41, N702);
xor XOR2_182 (N735, N45, N703);
xor XOR2_183 (N736, N49, N704);
xor XOR2_184 (N737, N53, N705);
xor XOR2_185 (N738, N57, N706);
xor XOR2_186 (N739, N61, N707);
xor XOR2_187 (N740, N65, N708);
xor XOR2_188 (N741, N69, N709);
xor XOR2_189 (N742, N73, N710);
xor XOR2_190 (N743, N77, N711);
xor XOR2_191 (N744, N81, N712);
xor XOR2_192 (N745, N85, N713);
xor XOR2_193 (N746, N89, N714);
xor XOR2_194 (N747, N93, N715);
xor XOR2_195 (N748, N97, N716);
xor XOR2_196 (N749, N101, N717);
xor XOR2_197 (N750, N105, N718);
xor XOR2_198 (N751, N109, N719);
xor XOR2_199 (N752, N113, N720);
xor XOR2_200 (N753, N117, N721);
xor XOR2_201 (N754, N121, N722);
xor XOR2_202 (N755, N125, N723);

endmodule
