`timescale 1ns / 1ps
// Verilog
// c432
// Ninputs 36
// Noutputs 7
// NtotalGates 160
// NOT1 40
// NAND2 64
// NOR2 19
// AND9 3
// XOR2 18
// NAND4 14
// AND8 1
// NAND3 1

module top (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
                  N430,N431,N432,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
        keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
                  keyinput125, keyinput126, keyinput127,
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
                  keyinput198, keyinput199,
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
        keyinput235);

  input keyinput200, keyinput201, keyinput202, keyinput203, keyinput204;
  input keyinput205, keyinput206, keyinput207, keyinput208, keyinput209;
  input keyinput210, keyinput211, keyinput212, keyinput213, keyinput214;
  input keyinput215, keyinput216, keyinput217, keyinput218, keyinput219;
  input keyinput220, keyinput221, keyinput222, keyinput223, keyinput224;
  input keyinput225, keyinput226, keyinput227, keyinput228, keyinput229;
  input keyinput230, keyinput231, keyinput232, keyinput233, keyinput234;
  input keyinput235;


  input keyinput128, keyinput129, keyinput130, keyinput131, keyinput132;
  input keyinput133, keyinput134, keyinput135, keyinput136, keyinput137;
  input keyinput138, keyinput139, keyinput140, keyinput141, keyinput142;
  input keyinput143, keyinput144, keyinput145, keyinput146, keyinput147;
  input keyinput148, keyinput149, keyinput150, keyinput151, keyinput152;
  input keyinput153, keyinput154, keyinput155, keyinput156, keyinput157;
  input keyinput158, keyinput159, keyinput160, keyinput161, keyinput162;
  input keyinput163, keyinput164, keyinput165, keyinput166, keyinput167;
  input keyinput168, keyinput169, keyinput170, keyinput171, keyinput172;
  input keyinput173, keyinput174, keyinput175, keyinput176, keyinput177;
  input keyinput178, keyinput179, keyinput180, keyinput181, keyinput182;
  input keyinput183, keyinput184, keyinput185, keyinput186, keyinput187;
  input keyinput188, keyinput189, keyinput190, keyinput191, keyinput192;
  input keyinput193, keyinput194, keyinput195, keyinput196, keyinput197;
  input keyinput198, keyinput199;

  wire KeyWire_0_1 , KeyWire_0_2;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31, keyinput32, keyinput33, keyinput34;
  input keyinput35, keyinput36, keyinput37, keyinput38, keyinput39;
  input keyinput40, keyinput41, keyinput42, keyinput43, keyinput44;
  input keyinput45, keyinput46, keyinput47, keyinput48, keyinput49;
  input keyinput50, keyinput51, keyinput52, keyinput53, keyinput54;
  input keyinput55, keyinput56, keyinput57, keyinput58, keyinput59;
  input keyinput60, keyinput61, keyinput62, keyinput63, keyinput64;
  input keyinput65, keyinput66, keyinput67, keyinput68, keyinput69;
  input keyinput70, keyinput71, keyinput72, keyinput73, keyinput74;
  input keyinput75, keyinput76, keyinput77, keyinput78, keyinput79;
  input keyinput80, keyinput81, keyinput82, keyinput83, keyinput84;
  input keyinput85, keyinput86, keyinput87, keyinput88, keyinput89;
  input keyinput90, keyinput91, keyinput92, keyinput93, keyinput94;
  input keyinput95, keyinput96, keyinput97, keyinput98, keyinput99;
  input keyinput100, keyinput101, keyinput102, keyinput103, keyinput104;
  input keyinput105, keyinput106, keyinput107, keyinput108, keyinput109;
  input keyinput110, keyinput111, keyinput112, keyinput113, keyinput114;
  input keyinput115, keyinput116, keyinput117, keyinput118, keyinput119;
  input keyinput120, keyinput121, keyinput122, keyinput123, keyinput124;
  input keyinput125, keyinput126, keyinput127;

  wire [0:127] keyinput_Wire_0;
  wire [0:66] KeyNOTWire_0;

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;

output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429;

  not NOT1_1 (keyinput_Wire_0[0], N1);
  xor keyGate_0_0(N118, keyinput0, keyinput_Wire_0[0]);
  not NOT1_2 (keyinput_Wire_0[1], N4);
  xor keyGate_0_1(KeyNOTWire_0[0], keyinput1, keyinput_Wire_0[1]);
  not KeyNOTGate_0_0(N119, KeyNOTWire_0[0]);
  not NOT1_3 (keyinput_Wire_0[2], N11);
  xor keyGate_0_2(KeyNOTWire_0[1], keyinput2, keyinput_Wire_0[2]);
  not KeyNOTGate_0_1(N122, KeyNOTWire_0[1]);
  not NOT1_4 (keyinput_Wire_0[3], N17);
  xnor keyGate_0_3(KeyNOTWire_0[2], keyinput3, keyinput_Wire_0[3]);
  not KeyNOTGate_0_2(N123, KeyNOTWire_0[2]);
  not NOT1_5 (keyinput_Wire_0[4], N24);
  xnor keyGate_0_4(KeyNOTWire_0[3], keyinput4, keyinput_Wire_0[4]);
  not KeyNOTGate_0_3(N126, KeyNOTWire_0[3]);
not NOT1_6 (N127, N30);
  not NOT1_7 (keyinput_Wire_0[5], N37);
  xor keyGate_0_5(N130, keyinput5, keyinput_Wire_0[5]);
not NOT1_8 (N131, N43);
  not NOT1_9 (keyinput_Wire_0[6], N50);
  xor keyGate_0_6(KeyNOTWire_0[4], keyinput6, keyinput_Wire_0[6]);
  not KeyNOTGate_0_4(N134, KeyNOTWire_0[4]);
  not NOT1_10 (keyinput_Wire_0[7], N56);
  xor keyGate_0_7(KeyNOTWire_0[5], keyinput7, keyinput_Wire_0[7]);
  not KeyNOTGate_0_5(N135, KeyNOTWire_0[5]);
not NOT1_11 (N138, N63);
  not NOT1_12 (keyinput_Wire_0[8], N69);
  xnor keyGate_0_8(KeyNOTWire_0[6], keyinput8, keyinput_Wire_0[8]);
  not KeyNOTGate_0_6(N139, KeyNOTWire_0[6]);
  not NOT1_13 (keyinput_Wire_0[9], N76);
  xor keyGate_0_9(N142, keyinput9, keyinput_Wire_0[9]);
not NOT1_14 (N143, N82);
  not NOT1_15 (keyinput_Wire_0[10], N89);
  xnor keyGate_0_10(N146, keyinput10, keyinput_Wire_0[10]);
not NOT1_16 (N147, N95);
  not NOT1_17 (keyinput_Wire_0[11], N102);
  xnor keyGate_0_11(N150, keyinput11, keyinput_Wire_0[11]);
  not NOT1_18 (keyinput_Wire_0[12], N108);
  xor keyGate_0_12(N151, keyinput12, keyinput_Wire_0[12]);
  nand NAND2_19 (keyinput_Wire_0[13], N118, N4);
  xor keyGate_0_13(N154, keyinput13, keyinput_Wire_0[13]);
  nor NOR2_20 (keyinput_Wire_0[14], N8, N119);
  xor keyGate_0_14(N157, keyinput14, keyinput_Wire_0[14]);
  nor NOR2_21 (keyinput_Wire_0[15], N14, N119);
  xnor keyGate_0_15(KeyNOTWire_0[7], keyinput15, keyinput_Wire_0[15]);
  not KeyNOTGate_0_7(N158, KeyNOTWire_0[7]);
nand NAND2_22 (N159, N122, N17);
  nand NAND2_23 (keyinput_Wire_0[16], N126, N30);
  xnor keyGate_0_16(KeyNOTWire_0[8], keyinput16, keyinput_Wire_0[16]);
  not KeyNOTGate_0_8(N162, KeyNOTWire_0[8]);
nand NAND2_24 (N165, N130, N43);
  nand NAND2_25 (keyinput_Wire_0[17], N134, N56);
  xor keyGate_0_17(N168, keyinput17, keyinput_Wire_0[17]);
  nand NAND2_26 (keyinput_Wire_0[18], N138, N69);
  xor keyGate_0_18(KeyNOTWire_0[9], keyinput18, keyinput_Wire_0[18]);
  not KeyNOTGate_0_9(N171, KeyNOTWire_0[9]);
nand NAND2_27 (N174, N142, N82);
  nand NAND2_28 (keyinput_Wire_0[19], N146, N95);
  xor keyGate_0_19(N177, keyinput19, keyinput_Wire_0[19]);
nand NAND2_29 (N180, N150, N108);
  nor NOR2_30 (keyinput_Wire_0[20], N21, N123);
  xor keyGate_0_20(N183, keyinput20, keyinput_Wire_0[20]);
  nor NOR2_31 (keyinput_Wire_0[21], N27, N123);
  xnor keyGate_0_21(KeyNOTWire_0[10], keyinput21, keyinput_Wire_0[21]);
  not KeyNOTGate_0_10(N184, KeyNOTWire_0[10]);
  nor NOR2_32 (keyinput_Wire_0[22], N34, N127);
  xor keyGate_0_22(N185, keyinput22, keyinput_Wire_0[22]);
  nor NOR2_33 (keyinput_Wire_0[23], N40, N127);
  xnor keyGate_0_23(N186, keyinput23, keyinput_Wire_0[23]);
  nor NOR2_34 (keyinput_Wire_0[24], N47, N131);
  xor keyGate_0_24(N187, keyinput24, keyinput_Wire_0[24]);
  nor NOR2_35 (keyinput_Wire_0[25], N53, N131);
  xor keyGate_0_25(KeyNOTWire_0[11], keyinput25, keyinput_Wire_0[25]);
  not KeyNOTGate_0_11(N188, KeyNOTWire_0[11]);
  nor NOR2_36 (keyinput_Wire_0[26], N60, N135);
  xor keyGate_0_26(KeyNOTWire_0[12], keyinput26, keyinput_Wire_0[26]);
  not KeyNOTGate_0_12(N189, KeyNOTWire_0[12]);
  nor NOR2_37 (keyinput_Wire_0[27], N66, N135);
  xnor keyGate_0_27(KeyNOTWire_0[13], keyinput27, keyinput_Wire_0[27]);
  not KeyNOTGate_0_13(N190, KeyNOTWire_0[13]);
  nor NOR2_38 (keyinput_Wire_0[28], N73, N139);
  xor keyGate_0_28(KeyNOTWire_0[14], keyinput28, keyinput_Wire_0[28]);
  not KeyNOTGate_0_14(N191, KeyNOTWire_0[14]);
  nor NOR2_39 (keyinput_Wire_0[29], N79, N139);
  xnor keyGate_0_29(N192, keyinput29, keyinput_Wire_0[29]);
  nor NOR2_40 (keyinput_Wire_0[30], N86, N143);
  xnor keyGate_0_30(KeyNOTWire_0[15], keyinput30, keyinput_Wire_0[30]);
  not KeyNOTGate_0_15(N193, KeyNOTWire_0[15]);
nor NOR2_41 (N194, N92, N143);
  nor NOR2_42 (keyinput_Wire_0[31], N99, N147);
  xnor keyGate_0_31(KeyNOTWire_0[16], keyinput31, keyinput_Wire_0[31]);
  not KeyNOTGate_0_16(N195, KeyNOTWire_0[16]);
  nor NOR2_43 (keyinput_Wire_0[32], N105, N147);
  xor keyGate_0_32(KeyNOTWire_0[17], keyinput32, keyinput_Wire_0[32]);
  not KeyNOTGate_0_17(N196, KeyNOTWire_0[17]);
  nor NOR2_44 (keyinput_Wire_0[33], N112, N151);
  xor keyGate_0_33(KeyNOTWire_0[18], keyinput33, keyinput_Wire_0[33]);
  not KeyNOTGate_0_18(N197, KeyNOTWire_0[18]);
nor NOR2_45 (N198, N115, N151);
  and AND9_46 (keyinput_Wire_0[34], N154, N159, N162, N165, N168, N171, N174, N177, N180);
  xor keyGate_0_34(N199, keyinput34, keyinput_Wire_0[34]);
  not NOT1_47 (keyinput_Wire_0[35], N199);
  xnor keyGate_0_35(N203, keyinput35, keyinput_Wire_0[35]);
not NOT1_48 (N213, N199);
not NOT1_49 (N223, N199);
xor XOR2_50 (N224, N203, N154);
  xor XOR2_51 (keyinput_Wire_0[36], N203, N159);
  xnor keyGate_0_36(KeyNOTWire_0[19], keyinput36, keyinput_Wire_0[36]);
  not KeyNOTGate_0_19(N227, KeyNOTWire_0[19]);
  xor XOR2_52 (keyinput_Wire_0[37], N203, N162);
  xor keyGate_0_37(KeyNOTWire_0[20], keyinput37, keyinput_Wire_0[37]);
  not KeyNOTGate_0_20(N230, KeyNOTWire_0[20]);
  xor XOR2_53 (keyinput_Wire_0[38], N203, N165);
  xnor keyGate_0_38(KeyNOTWire_0[21], keyinput38, keyinput_Wire_0[38]);
  not KeyNOTGate_0_21(N233, KeyNOTWire_0[21]);
  xor XOR2_54 (keyinput_Wire_0[39], N203, N168);
  xor keyGate_0_39(N236, keyinput39, keyinput_Wire_0[39]);
  xor XOR2_55 (keyinput_Wire_0[40], N203, N171);
  xor keyGate_0_40(KeyNOTWire_0[22], keyinput40, keyinput_Wire_0[40]);
  not KeyNOTGate_0_22(N239, KeyNOTWire_0[22]);
  nand NAND2_56 (keyinput_Wire_0[41], N1, N213);
  xnor keyGate_0_41(KeyNOTWire_0[23], keyinput41, keyinput_Wire_0[41]);
  not KeyNOTGate_0_23(N242, KeyNOTWire_0[23]);
xor XOR2_57 (N243, N203, N174);
  nand NAND2_58 (keyinput_Wire_0[42], N213, N11);
  xor keyGate_0_42(KeyNOTWire_0[24], keyinput42, keyinput_Wire_0[42]);
  not KeyNOTGate_0_24(N246, KeyNOTWire_0[24]);
  xor XOR2_59 (keyinput_Wire_0[43], N203, N177);
  xor keyGate_0_43(KeyNOTWire_0[25], keyinput43, keyinput_Wire_0[43]);
  not KeyNOTGate_0_25(N247, KeyNOTWire_0[25]);
  nand NAND2_60 (keyinput_Wire_0[44], N213, N24);
  xnor keyGate_0_44(N250, keyinput44, keyinput_Wire_0[44]);
  xor XOR2_61 (keyinput_Wire_0[45], N203, N180);
  xnor keyGate_0_45(N251, keyinput45, keyinput_Wire_0[45]);
nand NAND2_62 (N254, N213, N37);
nand NAND2_63 (N255, N213, N50);
nand NAND2_64 (N256, N213, N63);
  nand NAND2_65 (keyinput_Wire_0[46], N213, N76);
  xor keyGate_0_46(KeyNOTWire_0[26], keyinput46, keyinput_Wire_0[46]);
  not KeyNOTGate_0_26(N257, KeyNOTWire_0[26]);
  nand NAND2_66 (keyinput_Wire_0[47], N213, N89);
  xor keyGate_0_47(N258, keyinput47, keyinput_Wire_0[47]);
  nand NAND2_67 (keyinput_Wire_0[48], N213, N102);
  xor keyGate_0_48(N259, keyinput48, keyinput_Wire_0[48]);
nand NAND2_68 (N260, N224, N157);
  nand NAND2_69 (keyinput_Wire_0[49], N224, N158);
  xnor keyGate_0_49(N263, keyinput49, keyinput_Wire_0[49]);
  nand NAND2_70 (keyinput_Wire_0[50], N227, N183);
  xnor keyGate_0_50(KeyNOTWire_0[27], keyinput50, keyinput_Wire_0[50]);
  not KeyNOTGate_0_27(N264, KeyNOTWire_0[27]);
  nand NAND2_71 (keyinput_Wire_0[51], N230, N185);
  xnor keyGate_0_51(N267, keyinput51, keyinput_Wire_0[51]);
  nand NAND2_72 (keyinput_Wire_0[52], N233, N187);
  xnor keyGate_0_52(KeyNOTWire_0[28], keyinput52, keyinput_Wire_0[52]);
  not KeyNOTGate_0_28(N270, KeyNOTWire_0[28]);
nand NAND2_73 (N273, N236, N189);
  nand NAND2_74 (keyinput_Wire_0[53], N239, N191);
  xnor keyGate_0_53(KeyNOTWire_0[29], keyinput53, keyinput_Wire_0[53]);
  not KeyNOTGate_0_29(N276, KeyNOTWire_0[29]);
  nand NAND2_75 (keyinput_Wire_0[54], N243, N193);
  xnor keyGate_0_54(KeyNOTWire_0[30], keyinput54, keyinput_Wire_0[54]);
  not KeyNOTGate_0_30(N279, KeyNOTWire_0[30]);
  nand NAND2_76 (keyinput_Wire_0[55], N247, N195);
  xnor keyGate_0_55(N282, keyinput55, keyinput_Wire_0[55]);
  nand NAND2_77 (keyinput_Wire_0[56], N251, N197);
  xor keyGate_0_56(N285, keyinput56, keyinput_Wire_0[56]);
  nand NAND2_78 (keyinput_Wire_0[57], N227, N184);
  xor keyGate_0_57(N288, keyinput57, keyinput_Wire_0[57]);
  nand NAND2_79 (keyinput_Wire_0[58], N230, N186);
  xor keyGate_0_58(N289, keyinput58, keyinput_Wire_0[58]);
  nand NAND2_80 (keyinput_Wire_0[59], N233, N188);
  xnor keyGate_0_59(N290, keyinput59, keyinput_Wire_0[59]);
  nand NAND2_81 (keyinput_Wire_0[60], N236, N190);
  xor keyGate_0_60(N291, keyinput60, keyinput_Wire_0[60]);
nand NAND2_82 (N292, N239, N192);
  nand NAND2_83 (keyinput_Wire_0[61], N243, N194);
  xor keyGate_0_61(KeyNOTWire_0[31], keyinput61, keyinput_Wire_0[61]);
  not KeyNOTGate_0_31(N293, KeyNOTWire_0[31]);
  nand NAND2_84 (keyinput_Wire_0[62], N247, N196);
  xnor keyGate_0_62(KeyNOTWire_0[32], keyinput62, keyinput_Wire_0[62]);
  not KeyNOTGate_0_32(N294, KeyNOTWire_0[32]);
  nand NAND2_85 (keyinput_Wire_0[63], N251, N198);
  xor keyGate_0_63(KeyNOTWire_0[33], keyinput63, keyinput_Wire_0[63]);
  not KeyNOTGate_0_33(N295, KeyNOTWire_0[33]);
and AND9_86 (N296, N260, N264, N267, N270, N273, N276, N279, N282, N285);
  not NOT1_87 (keyinput_Wire_0[64], N263);
  xor keyGate_0_64(KeyNOTWire_0[34], keyinput64, keyinput_Wire_0[64]);
  not KeyNOTGate_0_34(N300, KeyNOTWire_0[34]);
  not NOT1_88 (keyinput_Wire_0[65], N288);
  xor keyGate_0_65(N301, keyinput65, keyinput_Wire_0[65]);
  not NOT1_89 (keyinput_Wire_0[66], N289);
  xor keyGate_0_66(KeyNOTWire_0[35], keyinput66, keyinput_Wire_0[66]);
  not KeyNOTGate_0_35(N302, KeyNOTWire_0[35]);
  not NOT1_90 (keyinput_Wire_0[67], N290);
  xor keyGate_0_67(KeyNOTWire_0[36], keyinput67, keyinput_Wire_0[67]);
  not KeyNOTGate_0_36(N303, KeyNOTWire_0[36]);
  not NOT1_91 (keyinput_Wire_0[68], N291);
  xnor keyGate_0_68(N304, keyinput68, keyinput_Wire_0[68]);
  not NOT1_92 (keyinput_Wire_0[69], N292);
  xor keyGate_0_69(N305, keyinput69, keyinput_Wire_0[69]);
  not NOT1_93 (keyinput_Wire_0[70], N293);
  xor keyGate_0_70(KeyNOTWire_0[37], keyinput70, keyinput_Wire_0[70]);
  not KeyNOTGate_0_37(N306, KeyNOTWire_0[37]);
  not NOT1_94 (keyinput_Wire_0[71], N294);
  xnor keyGate_0_71(N307, keyinput71, keyinput_Wire_0[71]);
  not NOT1_95 (keyinput_Wire_0[72], N295);
  xor keyGate_0_72(KeyNOTWire_0[38], keyinput72, keyinput_Wire_0[72]);
  not KeyNOTGate_0_38(N308, KeyNOTWire_0[38]);
  not NOT1_96 (keyinput_Wire_0[73], N296);
  xnor keyGate_0_73(N309, keyinput73, keyinput_Wire_0[73]);
  not NOT1_97 (keyinput_Wire_0[74], N296);
  xor keyGate_0_74(N319, keyinput74, keyinput_Wire_0[74]);
  not NOT1_98 (keyinput_Wire_0[75], N296);
  xor keyGate_0_75(N329, keyinput75, keyinput_Wire_0[75]);
  xor XOR2_99 (keyinput_Wire_0[76], N309, N260);
  xnor keyGate_0_76(KeyNOTWire_0[39], keyinput76, keyinput_Wire_0[76]);
  not KeyNOTGate_0_39(N330, KeyNOTWire_0[39]);
  xor XOR2_100 (keyinput_Wire_0[77], N309, N264);
  xor keyGate_0_77(N331, keyinput77, keyinput_Wire_0[77]);
  xor XOR2_101 (keyinput_Wire_0[78], N309, N267);
  xor keyGate_0_78(N332, keyinput78, keyinput_Wire_0[78]);
  xor XOR2_102 (keyinput_Wire_0[79], N309, N270);
  xnor keyGate_0_79(KeyNOTWire_0[40], keyinput79, keyinput_Wire_0[79]);
  not KeyNOTGate_0_40(N333, KeyNOTWire_0[40]);
  nand NAND2_103 (keyinput_Wire_0[80], N8, N319);
  xnor keyGate_0_80(N334, keyinput80, keyinput_Wire_0[80]);
  xor XOR2_104 (keyinput_Wire_0[81], N309, N273);
  xor keyGate_0_81(KeyNOTWire_0[41], keyinput81, keyinput_Wire_0[81]);
  not KeyNOTGate_0_41(N335, KeyNOTWire_0[41]);
  nand NAND2_105 (keyinput_Wire_0[82], N319, N21);
  xor keyGate_0_82(KeyNOTWire_0[42], keyinput82, keyinput_Wire_0[82]);
  not KeyNOTGate_0_42(N336, KeyNOTWire_0[42]);
  xor XOR2_106 (keyinput_Wire_0[83], N309, N276);
  xor keyGate_0_83(N337, keyinput83, keyinput_Wire_0[83]);
  nand NAND2_107 (keyinput_Wire_0[84], N319, N34);
  xnor keyGate_0_84(KeyNOTWire_0[43], keyinput84, keyinput_Wire_0[84]);
  not KeyNOTGate_0_43(N338, KeyNOTWire_0[43]);
  xor XOR2_108 (keyinput_Wire_0[85], N309, N279);
  xor keyGate_0_85(N339, keyinput85, keyinput_Wire_0[85]);
  nand NAND2_109 (keyinput_Wire_0[86], N319, N47);
  xnor keyGate_0_86(N340, keyinput86, keyinput_Wire_0[86]);
  xor XOR2_110 (keyinput_Wire_0[87], N309, N282);
  xnor keyGate_0_87(N341, keyinput87, keyinput_Wire_0[87]);
  nand NAND2_111 (keyinput_Wire_0[88], N319, N60);
  xnor keyGate_0_88(KeyNOTWire_0[44], keyinput88, keyinput_Wire_0[88]);
  not KeyNOTGate_0_44(N342, KeyNOTWire_0[44]);
  xor XOR2_112 (keyinput_Wire_0[89], N309, N285);
  xnor keyGate_0_89(KeyNOTWire_0[45], keyinput89, keyinput_Wire_0[89]);
  not KeyNOTGate_0_45(N343, KeyNOTWire_0[45]);
nand NAND2_113 (N344, N319, N73);
  nand NAND2_114 (keyinput_Wire_0[90], N319, N86);
  xnor keyGate_0_90(KeyNOTWire_0[46], keyinput90, keyinput_Wire_0[90]);
  not KeyNOTGate_0_46(N345, KeyNOTWire_0[46]);
  nand NAND2_115 (keyinput_Wire_0[91], N319, N99);
  xnor keyGate_0_91(KeyNOTWire_0[47], keyinput91, keyinput_Wire_0[91]);
  not KeyNOTGate_0_47(N346, KeyNOTWire_0[47]);
  nand NAND2_116 (keyinput_Wire_0[92], N319, N112);
  xor keyGate_0_92(KeyNOTWire_0[48], keyinput92, keyinput_Wire_0[92]);
  not KeyNOTGate_0_48(N347, KeyNOTWire_0[48]);
nand NAND2_117 (N348, N330, N300);
nand NAND2_118 (N349, N331, N301);
  nand NAND2_119 (keyinput_Wire_0[93], N332, N302);
  xor keyGate_0_93(KeyNOTWire_0[49], keyinput93, keyinput_Wire_0[93]);
  not KeyNOTGate_0_49(N350, KeyNOTWire_0[49]);
  nand NAND2_120 (keyinput_Wire_0[94], N333, N303);
  xnor keyGate_0_94(N351, keyinput94, keyinput_Wire_0[94]);
  nand NAND2_121 (keyinput_Wire_0[95], N335, N304);
  xnor keyGate_0_95(N352, keyinput95, keyinput_Wire_0[95]);
nand NAND2_122 (N353, N337, N305);
  nand NAND2_123 (keyinput_Wire_0[96], N339, N306);
  xor keyGate_0_96(N354, keyinput96, keyinput_Wire_0[96]);
  nand NAND2_124 (keyinput_Wire_0[97], N341, N307);
  xor keyGate_0_97(KeyNOTWire_0[50], keyinput97, keyinput_Wire_0[97]);
  not KeyNOTGate_0_50(N355, KeyNOTWire_0[50]);
  nand NAND2_125 (keyinput_Wire_0[98], N343, N308);
  xor keyGate_0_98(KeyNOTWire_0[51], keyinput98, keyinput_Wire_0[98]);
  not KeyNOTGate_0_51(N356, KeyNOTWire_0[51]);
  and AND9_126 (keyinput_Wire_0[99], N348, N349, N350, N351, N352, N353, N354, N355, N356);
  xor keyGate_0_99(N357, keyinput99, keyinput_Wire_0[99]);
  not NOT1_127 (keyinput_Wire_0[100], N357);
  xnor keyGate_0_100(N360, keyinput100, keyinput_Wire_0[100]);
not NOT1_128 (KeyWire_0_1, N357);
  xor flip_it (N370, KeyWire_0_1, KeyWire_0_2 );
nand NAND2_129 (N371, N14, N360);
nand NAND2_130 (N372, N360, N27);
  nand NAND2_131 (keyinput_Wire_0[101], N360, N40);
  xnor keyGate_0_101(KeyNOTWire_0[52], keyinput101, keyinput_Wire_0[101]);
  not KeyNOTGate_0_52(N373, KeyNOTWire_0[52]);
  nand NAND2_132 (keyinput_Wire_0[102], N360, N53);
  xnor keyGate_0_102(KeyNOTWire_0[53], keyinput102, keyinput_Wire_0[102]);
  not KeyNOTGate_0_53(N374, KeyNOTWire_0[53]);
  nand NAND2_133 (keyinput_Wire_0[103], N360, N66);
  xor keyGate_0_103(N375, keyinput103, keyinput_Wire_0[103]);
nand NAND2_134 (N376, N360, N79);
  nand NAND2_135 (keyinput_Wire_0[104], N360, N92);
  xnor keyGate_0_104(N377, keyinput104, keyinput_Wire_0[104]);
  nand NAND2_136 (keyinput_Wire_0[105], N360, N105);
  xnor keyGate_0_105(N378, keyinput105, keyinput_Wire_0[105]);
  nand NAND2_137 (keyinput_Wire_0[106], N360, N115);
  xor keyGate_0_106(N379, keyinput106, keyinput_Wire_0[106]);
  nand NAND4_138 (keyinput_Wire_0[107], N4, N242, N334, N371);
  xnor keyGate_0_107(KeyNOTWire_0[54], keyinput107, keyinput_Wire_0[107]);
  not KeyNOTGate_0_54(N380, KeyNOTWire_0[54]);
  nand NAND4_139 (keyinput_Wire_0[108], N246, N336, N372, N17);
  xnor keyGate_0_108(KeyNOTWire_0[55], keyinput108, keyinput_Wire_0[108]);
  not KeyNOTGate_0_55(N381, KeyNOTWire_0[55]);
  nand NAND4_140 (keyinput_Wire_0[109], N250, N338, N373, N30);
  xnor keyGate_0_109(KeyNOTWire_0[56], keyinput109, keyinput_Wire_0[109]);
  not KeyNOTGate_0_56(N386, KeyNOTWire_0[56]);
  nand NAND4_141 (keyinput_Wire_0[110], N254, N340, N374, N43);
  xnor keyGate_0_110(N393, keyinput110, keyinput_Wire_0[110]);
  nand NAND4_142 (keyinput_Wire_0[111], N255, N342, N375, N56);
  xnor keyGate_0_111(N399, keyinput111, keyinput_Wire_0[111]);
nand NAND4_143 (N404, N256, N344, N376, N69);
  nand NAND4_144 (keyinput_Wire_0[112], N257, N345, N377, N82);
  xor keyGate_0_112(KeyNOTWire_0[57], keyinput112, keyinput_Wire_0[112]);
  not KeyNOTGate_0_57(N407, KeyNOTWire_0[57]);
  nand NAND4_145 (keyinput_Wire_0[113], N258, N346, N378, N95);
  xor keyGate_0_113(KeyNOTWire_0[58], keyinput113, keyinput_Wire_0[113]);
  not KeyNOTGate_0_58(N411, KeyNOTWire_0[58]);
  nand NAND4_146 (keyinput_Wire_0[114], N259, N347, N379, N108);
  xor keyGate_0_114(N414, keyinput114, keyinput_Wire_0[114]);
  not NOT1_147 (keyinput_Wire_0[115], N380);
  xor keyGate_0_115(N415, keyinput115, keyinput_Wire_0[115]);
  and AND8_148 (keyinput_Wire_0[116], N381, N386, N393, N399, N404, N407, N411, N414);
  xnor keyGate_0_116(KeyNOTWire_0[59], keyinput116, keyinput_Wire_0[116]);
  not KeyNOTGate_0_59(N416, KeyNOTWire_0[59]);
  not NOT1_149 (keyinput_Wire_0[117], N393);
  xnor keyGate_0_117(KeyNOTWire_0[60], keyinput117, keyinput_Wire_0[117]);
  not KeyNOTGate_0_60(N417, KeyNOTWire_0[60]);
  not NOT1_150 (keyinput_Wire_0[118], N404);
  xor keyGate_0_118(KeyNOTWire_0[61], keyinput118, keyinput_Wire_0[118]);
  not KeyNOTGate_0_61(N418, KeyNOTWire_0[61]);
  not NOT1_151 (keyinput_Wire_0[119], N407);
  xnor keyGate_0_119(N419, keyinput119, keyinput_Wire_0[119]);
  not NOT1_152 (keyinput_Wire_0[120], N411);
  xnor keyGate_0_120(KeyNOTWire_0[62], keyinput120, keyinput_Wire_0[120]);
  not KeyNOTGate_0_62(N420, KeyNOTWire_0[62]);
  nor NOR2_153 (keyinput_Wire_0[121], N415, N416);
  xor keyGate_0_121(KeyNOTWire_0[63], keyinput121, keyinput_Wire_0[121]);
  not KeyNOTGate_0_63(N421, KeyNOTWire_0[63]);
  nand NAND2_154 (keyinput_Wire_0[122], N386, N417);
  xnor keyGate_0_122(N422, keyinput122, keyinput_Wire_0[122]);
  nand NAND4_155 (keyinput_Wire_0[123], N386, N393, N418, N399);
  xnor keyGate_0_123(N425, keyinput123, keyinput_Wire_0[123]);
  nand NAND3_156 (keyinput_Wire_0[124], N399, N393, N419);
  xor keyGate_0_124(KeyNOTWire_0[64], keyinput124, keyinput_Wire_0[124]);
  not KeyNOTGate_0_64(N428, KeyNOTWire_0[64]);
  nand NAND4_157 (keyinput_Wire_0[125], N386, N393, N407, N420);
  xor keyGate_0_125(N429, keyinput125, keyinput_Wire_0[125]);
  nand NAND4_158 (keyinput_Wire_0[126], N381, N386, N422, N399);
  xor keyGate_0_126(KeyNOTWire_0[65], keyinput126, keyinput_Wire_0[126]);
  not KeyNOTGate_0_65(N430, KeyNOTWire_0[65]);
  nand NAND4_159 (keyinput_Wire_0[127], N381, N386, N425, N428);
  xnor keyGate_0_127(KeyNOTWire_0[66], keyinput127, keyinput_Wire_0[127]);
  not KeyNOTGate_0_66(N431, KeyNOTWire_0[66]);
nand NAND4_160 (N432, N381, N422, N425, N429);

AntiSAT some_name( KeyWire_0_2, N17, N105, N4, N11, N63, N69, N79, N47, N73, N50, N24, N108, N92, N86, N82, N34, N43, N40, N21, N99, N89, N30, N115, N56, N27, N66, N60, N102, N112, N95, N8, N1, N53, N37, N14, N76, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
       keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
       keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
       keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
       keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
       keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
       keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
       keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
       keyinput235);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N17, N105, N4, N11, N63, N69, N79, N47, N73, N50, N24, N108, N92, N86, N82, N34, N43, N40, N21, N99, N89, N30, N115, N56, N27, N66, N60, N102, N112, N95, N8, N1, N53, N37, N14, N76, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199 ,
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
        keyinput235);

  input keyinput200, keyinput201, keyinput202, keyinput203, keyinput204;
  input keyinput205, keyinput206, keyinput207, keyinput208, keyinput209;
  input keyinput210, keyinput211, keyinput212, keyinput213, keyinput214;
  input keyinput215, keyinput216, keyinput217, keyinput218, keyinput219;
  input keyinput220, keyinput221, keyinput222, keyinput223, keyinput224;
  input keyinput225, keyinput226, keyinput227, keyinput228, keyinput229;
  input keyinput230, keyinput231, keyinput232, keyinput233, keyinput234;
  input keyinput235;

  wire [0:35] keyNTin_Wire_1;
  wire [0:13] KeyNOTWire_1;

  input N17, N105, N4, N11, N63, N69, N79, N47, N73, N50, N24, N108, N92, N86, N82, N34, N43, N40, N21, N99, N89, N30, N115, N56, N27, N66, N60, N102, N112, N95, N8, N1, N53, N37, N14, N76;
  input keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73 ;

  xnor KeyGate0 (newWire_0, N17, keyinput128);
  xnor KeyGate1 (keyNTin_Wire_1[0], N105, keyinput129);
  xor keyNTinGate_1_0(newWire_1, keyinput200, keyNTin_Wire_1[0]);
  xor  KeyGate2 (keyNTin_Wire_1[1], N4, keyinput130);
  xor keyNTinGate_1_1(newWire_2, keyinput201, keyNTin_Wire_1[1]);
  xor  KeyGate3 (newWire_3, N11, keyinput131);
  xnor KeyGate4 (keyNTin_Wire_1[2], N63, keyinput132);
  xnor keyNTinGate_1_2(KeyNOTWire_1[0], keyinput202, keyNTin_Wire_1[2]);
  not KeyNOTGate_1_0(newWire_4, KeyNOTWire_1[0]);
  xor  KeyGate5 (newWire_5, N69, keyinput133);
  xnor KeyGate6 (keyNTin_Wire_1[3], N79, keyinput134);
  xnor keyNTinGate_1_3(newWire_6, keyinput203, keyNTin_Wire_1[3]);
  xnor KeyGate7 (newWire_7, N47, keyinput135);
  xor  KeyGate8 (newWire_8, N73, keyinput136);
  xor  KeyGate9 (newWire_9, N50, keyinput137);
  xnor KeyGate10 (newWire_10, N24, keyinput138);
  xor  KeyGate11 (keyNTin_Wire_1[4], N108, keyinput139);
  xnor keyNTinGate_1_4(newWire_11, keyinput204, keyNTin_Wire_1[4]);
  xnor KeyGate12 (keyNTin_Wire_1[5], N92, keyinput140);
  xor keyNTinGate_1_5(newWire_12, keyinput205, keyNTin_Wire_1[5]);
  xnor KeyGate13 (keyNTin_Wire_1[6], N86, keyinput141);
  xnor keyNTinGate_1_6(newWire_13, keyinput206, keyNTin_Wire_1[6]);
  xnor KeyGate14 (newWire_14, N82, keyinput142);
  xnor KeyGate15 (newWire_15, N34, keyinput143);
  xnor KeyGate16 (newWire_16, N43, keyinput144);
  xnor KeyGate17 (keyNTin_Wire_1[7], N40, keyinput145);
  xor keyNTinGate_1_7(newWire_17, keyinput207, keyNTin_Wire_1[7]);
  xnor KeyGate18 (keyNTin_Wire_1[8], N21, keyinput146);
  xor keyNTinGate_1_8(newWire_18, keyinput208, keyNTin_Wire_1[8]);
  xor  KeyGate19 (keyNTin_Wire_1[9], N99, keyinput147);
  xor keyNTinGate_1_9(KeyNOTWire_1[1], keyinput209, keyNTin_Wire_1[9]);
  not KeyNOTGate_1_1(newWire_19, KeyNOTWire_1[1]);
  xor  KeyGate20 (newWire_20, N89, keyinput148);
  xnor KeyGate21 (keyNTin_Wire_1[10], N30, keyinput149);
  xor keyNTinGate_1_10(KeyNOTWire_1[2], keyinput210, keyNTin_Wire_1[10]);
  not KeyNOTGate_1_2(newWire_21, KeyNOTWire_1[2]);
  xnor KeyGate22 (newWire_22, N115, keyinput150);
  xor  KeyGate23 (keyNTin_Wire_1[11], N56, keyinput151);
  xor keyNTinGate_1_11(newWire_23, keyinput211, keyNTin_Wire_1[11]);
  xor  KeyGate24 (keyNTin_Wire_1[12], N27, keyinput152);
  xor keyNTinGate_1_12(newWire_24, keyinput212, keyNTin_Wire_1[12]);
  xor  KeyGate25 (keyNTin_Wire_1[13], N66, keyinput153);
  xnor keyNTinGate_1_13(newWire_25, keyinput213, keyNTin_Wire_1[13]);
  xor  KeyGate26 (newWire_26, N60, keyinput154);
  xnor KeyGate27 (keyNTin_Wire_1[14], N102, keyinput155);
  xnor keyNTinGate_1_14(KeyNOTWire_1[3], keyinput214, keyNTin_Wire_1[14]);
  not KeyNOTGate_1_3(newWire_27, KeyNOTWire_1[3]);
  xnor KeyGate28 (newWire_28, N112, keyinput156);
  xor  KeyGate29 (keyNTin_Wire_1[15], N95, keyinput157);
  xor keyNTinGate_1_15(newWire_29, keyinput215, keyNTin_Wire_1[15]);
  xor  KeyGate30 (keyNTin_Wire_1[16], N8, keyinput158);
  xor keyNTinGate_1_16(newWire_30, keyinput216, keyNTin_Wire_1[16]);
  xnor KeyGate31 (keyNTin_Wire_1[17], N1, keyinput159);
  xnor keyNTinGate_1_17(newWire_31, keyinput217, keyNTin_Wire_1[17]);
  xnor KeyGate32 (newWire_32, N53, keyinput160);
  xor  KeyGate33 (keyNTin_Wire_1[18], N37, keyinput161);
  xnor keyNTinGate_1_18(KeyNOTWire_1[4], keyinput218, keyNTin_Wire_1[18]);
  not KeyNOTGate_1_4(newWire_33, KeyNOTWire_1[4]);
  xor  KeyGate34 (newWire_34, N14, keyinput162);
  xor  KeyGate35 (newWire_35, N76, keyinput163);
  xnor KeyGate36 (newWire_36, N17, keyinput164);
  xnor KeyGate37 (keyNTin_Wire_1[19], N105, keyinput165);
  xnor keyNTinGate_1_19(newWire_37, keyinput219, keyNTin_Wire_1[19]);
  xor  KeyGate38 (newWire_38, N4, keyinput166);
  xnor KeyGate39 (newWire_39, N11, keyinput167);
  xnor KeyGate40 (newWire_40, N63, keyinput168);
  xnor KeyGate41 (keyNTin_Wire_1[20], N69, keyinput169);
  xor keyNTinGate_1_20(KeyNOTWire_1[5], keyinput220, keyNTin_Wire_1[20]);
  not KeyNOTGate_1_5(newWire_41, KeyNOTWire_1[5]);
  xnor KeyGate42 (newWire_42, N79, keyinput170);
  xnor KeyGate43 (newWire_43, N47, keyinput171);
  xnor KeyGate44 (newWire_44, N73, keyinput172);
  xor  KeyGate45 (newWire_45, N50, keyinput173);
  xor  KeyGate46 (keyNTin_Wire_1[21], N24, keyinput174);
  xor keyNTinGate_1_21(newWire_46, keyinput221, keyNTin_Wire_1[21]);
  xnor KeyGate47 (newWire_47, N108, keyinput175);
  xnor KeyGate48 (keyNTin_Wire_1[22], N92, keyinput176);
  xnor keyNTinGate_1_22(newWire_48, keyinput222, keyNTin_Wire_1[22]);
  xor  KeyGate49 (newWire_49, N86, keyinput177);
  xnor KeyGate50 (keyNTin_Wire_1[23], N82, keyinput178);
  xnor keyNTinGate_1_23(KeyNOTWire_1[6], keyinput223, keyNTin_Wire_1[23]);
  not KeyNOTGate_1_6(newWire_50, KeyNOTWire_1[6]);
  xnor KeyGate51 (keyNTin_Wire_1[24], N34, keyinput179);
  xor keyNTinGate_1_24(KeyNOTWire_1[7], keyinput224, keyNTin_Wire_1[24]);
  not KeyNOTGate_1_7(newWire_51, KeyNOTWire_1[7]);
  xnor KeyGate52 (newWire_52, N43, keyinput180);
  xor  KeyGate53 (keyNTin_Wire_1[25], N40, keyinput181);
  xor keyNTinGate_1_25(newWire_53, keyinput225, keyNTin_Wire_1[25]);
  xor  KeyGate54 (newWire_54, N21, keyinput182);
  xnor KeyGate55 (keyNTin_Wire_1[26], N99, keyinput183);
  xor keyNTinGate_1_26(newWire_55, keyinput226, keyNTin_Wire_1[26]);
  xor  KeyGate56 (newWire_56, N89, keyinput184);
  xnor KeyGate57 (keyNTin_Wire_1[27], N30, keyinput185);
  xor keyNTinGate_1_27(KeyNOTWire_1[8], keyinput227, keyNTin_Wire_1[27]);
  not KeyNOTGate_1_8(newWire_57, KeyNOTWire_1[8]);
  xnor KeyGate58 (newWire_58, N115, keyinput186);
  xnor KeyGate59 (newWire_59, N56, keyinput187);
  xnor KeyGate60 (keyNTin_Wire_1[28], N27, keyinput188);
  xor keyNTinGate_1_28(KeyNOTWire_1[9], keyinput228, keyNTin_Wire_1[28]);
  not KeyNOTGate_1_9(newWire_60, KeyNOTWire_1[9]);
  xnor KeyGate61 (newWire_61, N66, keyinput189);
  xnor KeyGate62 (newWire_62, N60, keyinput190);
  xor  KeyGate63 (keyNTin_Wire_1[29], N102, keyinput191);
  xnor keyNTinGate_1_29(KeyNOTWire_1[10], keyinput229, keyNTin_Wire_1[29]);
  not KeyNOTGate_1_10(newWire_63, KeyNOTWire_1[10]);
  xor  KeyGate64 (newWire_64, N112, keyinput192);
  xnor KeyGate65 (keyNTin_Wire_1[30], N95, keyinput193);
  xnor keyNTinGate_1_30(newWire_65, keyinput230, keyNTin_Wire_1[30]);
  xor  KeyGate66 (keyNTin_Wire_1[31], N8, keyinput194);
  xor keyNTinGate_1_31(KeyNOTWire_1[11], keyinput231, keyNTin_Wire_1[31]);
  not KeyNOTGate_1_11(newWire_66, KeyNOTWire_1[11]);
  xnor KeyGate67 (keyNTin_Wire_1[32], N1, keyinput195);
  xnor keyNTinGate_1_32(newWire_67, keyinput232, keyNTin_Wire_1[32]);
  xnor KeyGate68 (keyNTin_Wire_1[33], N53, keyinput196);
  xor keyNTinGate_1_33(KeyNOTWire_1[12], keyinput233, keyNTin_Wire_1[33]);
  not KeyNOTGate_1_12(newWire_68, KeyNOTWire_1[12]);
  xnor KeyGate69 (newWire_69, N37, keyinput197);
  xor  KeyGate70 (newWire_70, N14, keyinput198);
  xnor KeyGate71 (newWire_71, N76, keyinput199);
  and some_function (keyNTin_Wire_1[34], newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35 );
  xor keyNTinGate_1_34(KeyNOTWire_1[13], keyinput234, keyNTin_Wire_1[34]);
  not KeyNOTGate_1_13(newWire_72, KeyNOTWire_1[13]);
  nand compl_function (keyNTin_Wire_1[35], newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71);
  xnor keyNTinGate_1_35(newWire_73, keyinput235, keyNTin_Wire_1[35]);
  and finalAND (KeyWire_0_2, newWire_72, newWire_73);

endmodule /* AntiSAT */
