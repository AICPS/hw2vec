`timescale 1ns / 1ps
// Verilog
// c499
// Ninputs 41
// Noutputs 32
// NtotalGates 202
// XOR2 104
// AND2 40
// NOT1 40
// AND4 8
// OR4 2
// AND5 8

module top (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
                  N753,N754,N755,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
        keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
                  keyinput125, keyinput126, keyinput127,
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202,
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207,
                  keyinput208, keyinput209,
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
        keyinput250);

  input keyinput210, keyinput211, keyinput212, keyinput213, keyinput214;
  input keyinput215, keyinput216, keyinput217, keyinput218, keyinput219;
  input keyinput220, keyinput221, keyinput222, keyinput223, keyinput224;
  input keyinput225, keyinput226, keyinput227, keyinput228, keyinput229;
  input keyinput230, keyinput231, keyinput232, keyinput233, keyinput234;
  input keyinput235, keyinput236, keyinput237, keyinput238, keyinput239;
  input keyinput240, keyinput241, keyinput242, keyinput243, keyinput244;
  input keyinput245, keyinput246, keyinput247, keyinput248, keyinput249;
  input keyinput250;


  input keyinput128, keyinput129, keyinput130, keyinput131, keyinput132;
  input keyinput133, keyinput134, keyinput135, keyinput136, keyinput137;
  input keyinput138, keyinput139, keyinput140, keyinput141, keyinput142;
  input keyinput143, keyinput144, keyinput145, keyinput146, keyinput147;
  input keyinput148, keyinput149, keyinput150, keyinput151, keyinput152;
  input keyinput153, keyinput154, keyinput155, keyinput156, keyinput157;
  input keyinput158, keyinput159, keyinput160, keyinput161, keyinput162;
  input keyinput163, keyinput164, keyinput165, keyinput166, keyinput167;
  input keyinput168, keyinput169, keyinput170, keyinput171, keyinput172;
  input keyinput173, keyinput174, keyinput175, keyinput176, keyinput177;
  input keyinput178, keyinput179, keyinput180, keyinput181, keyinput182;
  input keyinput183, keyinput184, keyinput185, keyinput186, keyinput187;
  input keyinput188, keyinput189, keyinput190, keyinput191, keyinput192;
  input keyinput193, keyinput194, keyinput195, keyinput196, keyinput197;
  input keyinput198, keyinput199, keyinput200, keyinput201, keyinput202;
  input keyinput203, keyinput204, keyinput205, keyinput206, keyinput207;
  input keyinput208, keyinput209;

  wire KeyWire_0_1 , KeyWire_0_2;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31, keyinput32, keyinput33, keyinput34;
  input keyinput35, keyinput36, keyinput37, keyinput38, keyinput39;
  input keyinput40, keyinput41, keyinput42, keyinput43, keyinput44;
  input keyinput45, keyinput46, keyinput47, keyinput48, keyinput49;
  input keyinput50, keyinput51, keyinput52, keyinput53, keyinput54;
  input keyinput55, keyinput56, keyinput57, keyinput58, keyinput59;
  input keyinput60, keyinput61, keyinput62, keyinput63, keyinput64;
  input keyinput65, keyinput66, keyinput67, keyinput68, keyinput69;
  input keyinput70, keyinput71, keyinput72, keyinput73, keyinput74;
  input keyinput75, keyinput76, keyinput77, keyinput78, keyinput79;
  input keyinput80, keyinput81, keyinput82, keyinput83, keyinput84;
  input keyinput85, keyinput86, keyinput87, keyinput88, keyinput89;
  input keyinput90, keyinput91, keyinput92, keyinput93, keyinput94;
  input keyinput95, keyinput96, keyinput97, keyinput98, keyinput99;
  input keyinput100, keyinput101, keyinput102, keyinput103, keyinput104;
  input keyinput105, keyinput106, keyinput107, keyinput108, keyinput109;
  input keyinput110, keyinput111, keyinput112, keyinput113, keyinput114;
  input keyinput115, keyinput116, keyinput117, keyinput118, keyinput119;
  input keyinput120, keyinput121, keyinput122, keyinput123, keyinput124;
  input keyinput125, keyinput126, keyinput127;

  wire [0:127] keyinput_Wire_0;
  wire [0:70] KeyNOTWire_0;

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;

output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723;

xor XOR2_1 (N250, N1, N5);
  xor XOR2_2 (keyinput_Wire_0[0], N9, N13);
  xnor keyGate_0_0(KeyNOTWire_0[0], keyinput0, keyinput_Wire_0[0]);
  not KeyNOTGate_0_0(N251, KeyNOTWire_0[0]);
xor XOR2_3 (N252, N17, N21);
  xor XOR2_4 (keyinput_Wire_0[1], N25, N29);
  xnor keyGate_0_1(KeyNOTWire_0[1], keyinput1, keyinput_Wire_0[1]);
  not KeyNOTGate_0_1(N253, KeyNOTWire_0[1]);
xor XOR2_5 (N254, N33, N37);
xor XOR2_6 (N255, N41, N45);
  xor XOR2_7 (keyinput_Wire_0[2], N49, N53);
  xor keyGate_0_2(KeyNOTWire_0[2], keyinput2, keyinput_Wire_0[2]);
  not KeyNOTGate_0_2(N256, KeyNOTWire_0[2]);
xor XOR2_8 (N257, N57, N61);
  xor XOR2_9 (keyinput_Wire_0[3], N65, N69);
  xnor keyGate_0_3(KeyNOTWire_0[3], keyinput3, keyinput_Wire_0[3]);
  not KeyNOTGate_0_3(N258, KeyNOTWire_0[3]);
  xor XOR2_10 (keyinput_Wire_0[4], N73, N77);
  xnor keyGate_0_4(KeyNOTWire_0[4], keyinput4, keyinput_Wire_0[4]);
  not KeyNOTGate_0_4(N259, KeyNOTWire_0[4]);
  xor XOR2_11 (keyinput_Wire_0[5], N81, N85);
  xor keyGate_0_5(KeyNOTWire_0[5], keyinput5, keyinput_Wire_0[5]);
  not KeyNOTGate_0_5(N260, KeyNOTWire_0[5]);
  xor XOR2_12 (keyinput_Wire_0[6], N89, N93);
  xnor keyGate_0_6(N261, keyinput6, keyinput_Wire_0[6]);
  xor XOR2_13 (keyinput_Wire_0[7], N97, N101);
  xor keyGate_0_7(N262, keyinput7, keyinput_Wire_0[7]);
  xor XOR2_14 (keyinput_Wire_0[8], N105, N109);
  xnor keyGate_0_8(N263, keyinput8, keyinput_Wire_0[8]);
  xor XOR2_15 (keyinput_Wire_0[9], N113, N117);
  xnor keyGate_0_9(N264, keyinput9, keyinput_Wire_0[9]);
  xor XOR2_16 (keyinput_Wire_0[10], N121, N125);
  xor keyGate_0_10(KeyNOTWire_0[6], keyinput10, keyinput_Wire_0[10]);
  not KeyNOTGate_0_6(N265, KeyNOTWire_0[6]);
  and AND2_17 (keyinput_Wire_0[11], N129, N137);
  xnor keyGate_0_11(KeyNOTWire_0[7], keyinput11, keyinput_Wire_0[11]);
  not KeyNOTGate_0_7(N266, KeyNOTWire_0[7]);
  and AND2_18 (keyinput_Wire_0[12], N130, N137);
  xnor keyGate_0_12(KeyNOTWire_0[8], keyinput12, keyinput_Wire_0[12]);
  not KeyNOTGate_0_8(N267, KeyNOTWire_0[8]);
and AND2_19 (N268, N131, N137);
  and AND2_20 (keyinput_Wire_0[13], N132, N137);
  xnor keyGate_0_13(KeyNOTWire_0[9], keyinput13, keyinput_Wire_0[13]);
  not KeyNOTGate_0_9(N269, KeyNOTWire_0[9]);
  and AND2_21 (keyinput_Wire_0[14], N133, N137);
  xor keyGate_0_14(KeyNOTWire_0[10], keyinput14, keyinput_Wire_0[14]);
  not KeyNOTGate_0_10(N270, KeyNOTWire_0[10]);
  and AND2_22 (keyinput_Wire_0[15], N134, N137);
  xor keyGate_0_15(N271, keyinput15, keyinput_Wire_0[15]);
  and AND2_23 (keyinput_Wire_0[16], N135, N137);
  xor keyGate_0_16(KeyNOTWire_0[11], keyinput16, keyinput_Wire_0[16]);
  not KeyNOTGate_0_11(N272, KeyNOTWire_0[11]);
  and AND2_24 (keyinput_Wire_0[17], N136, N137);
  xnor keyGate_0_17(N273, keyinput17, keyinput_Wire_0[17]);
xor XOR2_25 (N274, N1, N17);
xor XOR2_26 (N275, N33, N49);
xor XOR2_27 (N276, N5, N21);
  xor XOR2_28 (keyinput_Wire_0[18], N37, N53);
  xnor keyGate_0_18(N277, keyinput18, keyinput_Wire_0[18]);
xor XOR2_29 (N278, N9, N25);
  xor XOR2_30 (keyinput_Wire_0[19], N41, N57);
  xor keyGate_0_19(KeyNOTWire_0[12], keyinput19, keyinput_Wire_0[19]);
  not KeyNOTGate_0_12(N279, KeyNOTWire_0[12]);
  xor XOR2_31 (keyinput_Wire_0[20], N13, N29);
  xor keyGate_0_20(KeyNOTWire_0[13], keyinput20, keyinput_Wire_0[20]);
  not KeyNOTGate_0_13(N280, KeyNOTWire_0[13]);
xor XOR2_32 (N281, N45, N61);
  xor XOR2_33 (keyinput_Wire_0[21], N65, N81);
  xnor keyGate_0_21(N282, keyinput21, keyinput_Wire_0[21]);
  xor XOR2_34 (keyinput_Wire_0[22], N97, N113);
  xor keyGate_0_22(KeyNOTWire_0[14], keyinput22, keyinput_Wire_0[22]);
  not KeyNOTGate_0_14(N283, KeyNOTWire_0[14]);
  xor XOR2_35 (keyinput_Wire_0[23], N69, N85);
  xor keyGate_0_23(KeyNOTWire_0[15], keyinput23, keyinput_Wire_0[23]);
  not KeyNOTGate_0_15(N284, KeyNOTWire_0[15]);
xor XOR2_36 (N285, N101, N117);
  xor XOR2_37 (keyinput_Wire_0[24], N73, N89);
  xor keyGate_0_24(N286, keyinput24, keyinput_Wire_0[24]);
  xor XOR2_38 (keyinput_Wire_0[25], N105, N121);
  xnor keyGate_0_25(N287, keyinput25, keyinput_Wire_0[25]);
xor XOR2_39 (N288, N77, N93);
  xor XOR2_40 (keyinput_Wire_0[26], N109, N125);
  xnor keyGate_0_26(KeyNOTWire_0[16], keyinput26, keyinput_Wire_0[26]);
  not KeyNOTGate_0_16(N289, KeyNOTWire_0[16]);
  xor XOR2_41 (keyinput_Wire_0[27], N250, N251);
  xor keyGate_0_27(KeyNOTWire_0[17], keyinput27, keyinput_Wire_0[27]);
  not KeyNOTGate_0_17(N290, KeyNOTWire_0[17]);
  xor XOR2_42 (keyinput_Wire_0[28], N252, N253);
  xnor keyGate_0_28(KeyNOTWire_0[18], keyinput28, keyinput_Wire_0[28]);
  not KeyNOTGate_0_18(N293, KeyNOTWire_0[18]);
  xor XOR2_43 (keyinput_Wire_0[29], N254, N255);
  xnor keyGate_0_29(N296, keyinput29, keyinput_Wire_0[29]);
xor XOR2_44 (N299, N256, N257);
  xor XOR2_45 (keyinput_Wire_0[30], N258, N259);
  xor keyGate_0_30(N302, keyinput30, keyinput_Wire_0[30]);
  xor XOR2_46 (keyinput_Wire_0[31], N260, N261);
  xnor keyGate_0_31(N305, keyinput31, keyinput_Wire_0[31]);
  xor XOR2_47 (keyinput_Wire_0[32], N262, N263);
  xnor keyGate_0_32(N308, keyinput32, keyinput_Wire_0[32]);
  xor XOR2_48 (keyinput_Wire_0[33], N264, N265);
  xor keyGate_0_33(N311, keyinput33, keyinput_Wire_0[33]);
xor XOR2_49 (N314, N274, N275);
  xor XOR2_50 (keyinput_Wire_0[34], N276, N277);
  xnor keyGate_0_34(N315, keyinput34, keyinput_Wire_0[34]);
  xor XOR2_51 (keyinput_Wire_0[35], N278, N279);
  xnor keyGate_0_35(KeyNOTWire_0[19], keyinput35, keyinput_Wire_0[35]);
  not KeyNOTGate_0_19(N316, KeyNOTWire_0[19]);
  xor XOR2_52 (keyinput_Wire_0[36], N280, N281);
  xnor keyGate_0_36(KeyNOTWire_0[20], keyinput36, keyinput_Wire_0[36]);
  not KeyNOTGate_0_20(N317, KeyNOTWire_0[20]);
  xor XOR2_53 (keyinput_Wire_0[37], N282, N283);
  xor keyGate_0_37(KeyNOTWire_0[21], keyinput37, keyinput_Wire_0[37]);
  not KeyNOTGate_0_21(N318, KeyNOTWire_0[21]);
  xor XOR2_54 (keyinput_Wire_0[38], N284, N285);
  xnor keyGate_0_38(N319, keyinput38, keyinput_Wire_0[38]);
  xor XOR2_55 (keyinput_Wire_0[39], N286, N287);
  xor keyGate_0_39(N320, keyinput39, keyinput_Wire_0[39]);
  xor XOR2_56 (keyinput_Wire_0[40], N288, N289);
  xor keyGate_0_40(KeyNOTWire_0[22], keyinput40, keyinput_Wire_0[40]);
  not KeyNOTGate_0_22(N321, KeyNOTWire_0[22]);
xor XOR2_57 (N338, N290, N293);
  xor XOR2_58 (keyinput_Wire_0[41], N296, N299);
  xor keyGate_0_41(N339, keyinput41, keyinput_Wire_0[41]);
  xor XOR2_59 (keyinput_Wire_0[42], N290, N296);
  xor keyGate_0_42(KeyNOTWire_0[23], keyinput42, keyinput_Wire_0[42]);
  not KeyNOTGate_0_23(N340, KeyNOTWire_0[23]);
  xor XOR2_60 (keyinput_Wire_0[43], N293, N299);
  xor keyGate_0_43(KeyNOTWire_0[24], keyinput43, keyinput_Wire_0[43]);
  not KeyNOTGate_0_24(N341, KeyNOTWire_0[24]);
  xor XOR2_61 (keyinput_Wire_0[44], N302, N305);
  xor keyGate_0_44(KeyNOTWire_0[25], keyinput44, keyinput_Wire_0[44]);
  not KeyNOTGate_0_25(N342, KeyNOTWire_0[25]);
  xor XOR2_62 (keyinput_Wire_0[45], N308, N311);
  xnor keyGate_0_45(N343, keyinput45, keyinput_Wire_0[45]);
  xor XOR2_63 (keyinput_Wire_0[46], N302, N308);
  xor keyGate_0_46(KeyNOTWire_0[26], keyinput46, keyinput_Wire_0[46]);
  not KeyNOTGate_0_26(N344, KeyNOTWire_0[26]);
  xor XOR2_64 (keyinput_Wire_0[47], N305, N311);
  xor keyGate_0_47(KeyNOTWire_0[27], keyinput47, keyinput_Wire_0[47]);
  not KeyNOTGate_0_27(N345, KeyNOTWire_0[27]);
  xor XOR2_65 (keyinput_Wire_0[48], N266, N342);
  xor keyGate_0_48(KeyNOTWire_0[28], keyinput48, keyinput_Wire_0[48]);
  not KeyNOTGate_0_28(N346, KeyNOTWire_0[28]);
  xor XOR2_66 (keyinput_Wire_0[49], N267, N343);
  xnor keyGate_0_49(N347, keyinput49, keyinput_Wire_0[49]);
  xor XOR2_67 (keyinput_Wire_0[50], N268, N344);
  xnor keyGate_0_50(KeyNOTWire_0[29], keyinput50, keyinput_Wire_0[50]);
  not KeyNOTGate_0_29(N348, KeyNOTWire_0[29]);
  xor XOR2_68 (keyinput_Wire_0[51], N269, N345);
  xor keyGate_0_51(N349, keyinput51, keyinput_Wire_0[51]);
  xor XOR2_69 (keyinput_Wire_0[52], N270, N338);
  xnor keyGate_0_52(N350, keyinput52, keyinput_Wire_0[52]);
  xor XOR2_70 (keyinput_Wire_0[53], N271, N339);
  xnor keyGate_0_53(KeyNOTWire_0[30], keyinput53, keyinput_Wire_0[53]);
  not KeyNOTGate_0_30(N351, KeyNOTWire_0[30]);
  xor XOR2_71 (keyinput_Wire_0[54], N272, N340);
  xor keyGate_0_54(KeyNOTWire_0[31], keyinput54, keyinput_Wire_0[54]);
  not KeyNOTGate_0_31(N352, KeyNOTWire_0[31]);
xor XOR2_72 (N353, N273, N341);
xor XOR2_73 (N354, N314, N346);
xor XOR2_74 (N367, N315, N347);
  xor XOR2_75 (keyinput_Wire_0[55], N316, N348);
  xor keyGate_0_55(N380, keyinput55, keyinput_Wire_0[55]);
xor XOR2_76 (N393, N317, N349);
xor XOR2_77 (N406, N318, N350);
  xor XOR2_78 (keyinput_Wire_0[56], N319, N351);
  xnor keyGate_0_56(KeyNOTWire_0[32], keyinput56, keyinput_Wire_0[56]);
  not KeyNOTGate_0_32(N419, KeyNOTWire_0[32]);
xor XOR2_79 (N432, N320, N352);
xor XOR2_80 (N445, N321, N353);
  not NOT1_81 (keyinput_Wire_0[57], N354);
  xnor keyGate_0_57(KeyNOTWire_0[33], keyinput57, keyinput_Wire_0[57]);
  not KeyNOTGate_0_33(N554, KeyNOTWire_0[33]);
  not NOT1_82 (keyinput_Wire_0[58], N367);
  xnor keyGate_0_58(N555, keyinput58, keyinput_Wire_0[58]);
not NOT1_83 (N556, N380);
not NOT1_84 (N557, N354);
not NOT1_85 (N558, N367);
  not NOT1_86 (keyinput_Wire_0[59], N393);
  xor keyGate_0_59(KeyNOTWire_0[34], keyinput59, keyinput_Wire_0[59]);
  not KeyNOTGate_0_34(N559, KeyNOTWire_0[34]);
not NOT1_87 (N560, N354);
  not NOT1_88 (keyinput_Wire_0[60], N380);
  xor keyGate_0_60(KeyNOTWire_0[35], keyinput60, keyinput_Wire_0[60]);
  not KeyNOTGate_0_35(N561, KeyNOTWire_0[35]);
  not NOT1_89 (keyinput_Wire_0[61], N393);
  xnor keyGate_0_61(KeyNOTWire_0[36], keyinput61, keyinput_Wire_0[61]);
  not KeyNOTGate_0_36(N562, KeyNOTWire_0[36]);
not NOT1_90 (N563, N367);
  not NOT1_91 (keyinput_Wire_0[62], N380);
  xnor keyGate_0_62(N564, keyinput62, keyinput_Wire_0[62]);
  not NOT1_92 (keyinput_Wire_0[63], N393);
  xnor keyGate_0_63(N565, keyinput63, keyinput_Wire_0[63]);
not NOT1_93 (N566, N419);
not NOT1_94 (N567, N445);
  not NOT1_95 (keyinput_Wire_0[64], N419);
  xor keyGate_0_64(KeyNOTWire_0[37], keyinput64, keyinput_Wire_0[64]);
  not KeyNOTGate_0_37(N568, KeyNOTWire_0[37]);
  not NOT1_96 (keyinput_Wire_0[65], N432);
  xnor keyGate_0_65(KeyNOTWire_0[38], keyinput65, keyinput_Wire_0[65]);
  not KeyNOTGate_0_38(N569, KeyNOTWire_0[38]);
  not NOT1_97 (keyinput_Wire_0[66], N406);
  xnor keyGate_0_66(KeyNOTWire_0[39], keyinput66, keyinput_Wire_0[66]);
  not KeyNOTGate_0_39(N570, KeyNOTWire_0[39]);
  not NOT1_98 (keyinput_Wire_0[67], N445);
  xor keyGate_0_67(N571, keyinput67, keyinput_Wire_0[67]);
not NOT1_99 (N572, N406);
  not NOT1_100 (keyinput_Wire_0[68], N432);
  xnor keyGate_0_68(KeyNOTWire_0[40], keyinput68, keyinput_Wire_0[68]);
  not KeyNOTGate_0_40(N573, KeyNOTWire_0[40]);
  not NOT1_101 (keyinput_Wire_0[69], N406);
  xor keyGate_0_69(N574, keyinput69, keyinput_Wire_0[69]);
  not NOT1_102 (keyinput_Wire_0[70], N419);
  xor keyGate_0_70(N575, keyinput70, keyinput_Wire_0[70]);
not NOT1_103 (N576, N432);
not NOT1_104 (N577, N406);
  not NOT1_105 (keyinput_Wire_0[71], N419);
  xor keyGate_0_71(KeyNOTWire_0[41], keyinput71, keyinput_Wire_0[71]);
  not KeyNOTGate_0_41(N578, KeyNOTWire_0[41]);
not NOT1_106 (N579, N445);
  not NOT1_107 (keyinput_Wire_0[72], N406);
  xnor keyGate_0_72(KeyNOTWire_0[42], keyinput72, keyinput_Wire_0[72]);
  not KeyNOTGate_0_42(N580, KeyNOTWire_0[42]);
not NOT1_108 (N581, N432);
  not NOT1_109 (keyinput_Wire_0[73], N445);
  xor keyGate_0_73(N582, keyinput73, keyinput_Wire_0[73]);
  not NOT1_110 (keyinput_Wire_0[74], N419);
  xor keyGate_0_74(N583, keyinput74, keyinput_Wire_0[74]);
  not NOT1_111 (keyinput_Wire_0[75], N432);
  xnor keyGate_0_75(N584, keyinput75, keyinput_Wire_0[75]);
not NOT1_112 (N585, N445);
  not NOT1_113 (keyinput_Wire_0[76], N367);
  xnor keyGate_0_76(KeyNOTWire_0[43], keyinput76, keyinput_Wire_0[76]);
  not KeyNOTGate_0_43(N586, KeyNOTWire_0[43]);
  not NOT1_114 (keyinput_Wire_0[77], N393);
  xnor keyGate_0_77(KeyNOTWire_0[44], keyinput77, keyinput_Wire_0[77]);
  not KeyNOTGate_0_44(N587, KeyNOTWire_0[44]);
not NOT1_115 (N588, N367);
  not NOT1_116 (keyinput_Wire_0[78], N380);
  xor keyGate_0_78(N589, keyinput78, keyinput_Wire_0[78]);
  not NOT1_117 (keyinput_Wire_0[79], N354);
  xnor keyGate_0_79(N590, keyinput79, keyinput_Wire_0[79]);
not NOT1_118 (N591, N393);
not NOT1_119 (N592, N354);
not NOT1_120 (N593, N380);
  and AND4_121 (keyinput_Wire_0[80], N554, N555, N556, N393);
  xor keyGate_0_80(KeyNOTWire_0[45], keyinput80, keyinput_Wire_0[80]);
  not KeyNOTGate_0_45(N594, KeyNOTWire_0[45]);
  and AND4_122 (keyinput_Wire_0[81], N557, N558, N380, N559);
  xnor keyGate_0_81(KeyNOTWire_0[46], keyinput81, keyinput_Wire_0[81]);
  not KeyNOTGate_0_46(N595, KeyNOTWire_0[46]);
  and AND4_123 (keyinput_Wire_0[82], N560, N367, N561, N562);
  xor keyGate_0_82(N596, keyinput82, keyinput_Wire_0[82]);
  and AND4_124 (keyinput_Wire_0[83], N354, N563, N564, N565);
  xor keyGate_0_83(N597, keyinput83, keyinput_Wire_0[83]);
  and AND4_125 (keyinput_Wire_0[84], N574, N575, N576, N445);
  xnor keyGate_0_84(KeyNOTWire_0[47], keyinput84, keyinput_Wire_0[84]);
  not KeyNOTGate_0_47(N598, KeyNOTWire_0[47]);
and AND4_126 (N599, N577, N578, N432, N579);
and AND4_127 (N600, N580, N419, N581, N582);
  and AND4_128 (keyinput_Wire_0[85], N406, N583, N584, N585);
  xor keyGate_0_85(KeyNOTWire_0[48], keyinput85, keyinput_Wire_0[85]);
  not KeyNOTGate_0_48(N601, KeyNOTWire_0[48]);
  or OR4_129 (keyinput_Wire_0[86], N594, N595, N596, N597);
  xnor keyGate_0_86(KeyNOTWire_0[49], keyinput86, keyinput_Wire_0[86]);
  not KeyNOTGate_0_49(N602, KeyNOTWire_0[49]);
  or OR4_130 (keyinput_Wire_0[87], N598, N599, N600, N601);
  xor keyGate_0_87(KeyNOTWire_0[50], keyinput87, keyinput_Wire_0[87]);
  not KeyNOTGate_0_50(N607, KeyNOTWire_0[50]);
  and AND5_131 (keyinput_Wire_0[88], N406, N566, N432, N567, N602);
  xor keyGate_0_88(KeyNOTWire_0[51], keyinput88, keyinput_Wire_0[88]);
  not KeyNOTGate_0_51(N620, KeyNOTWire_0[51]);
  and AND5_132 (keyinput_Wire_0[89], N406, N568, N569, N445, N602);
  xnor keyGate_0_89(KeyNOTWire_0[52], keyinput89, keyinput_Wire_0[89]);
  not KeyNOTGate_0_52(N625, KeyNOTWire_0[52]);
and AND5_133 (N630, N570, N419, N432, N571, N602);
and AND5_134 (N635, N572, N419, N573, N445, N602);
  and AND5_135 (keyinput_Wire_0[90], N354, N586, N380, N587, N607);
  xnor keyGate_0_90(KeyNOTWire_0[53], keyinput90, keyinput_Wire_0[90]);
  not KeyNOTGate_0_53(N640, KeyNOTWire_0[53]);
and AND5_136 (N645, N354, N588, N589, N393, N607);
  and AND5_137 (keyinput_Wire_0[91], N590, N367, N380, N591, N607);
  xnor keyGate_0_91(N650, keyinput91, keyinput_Wire_0[91]);
and AND5_138 (N655, N592, N367, N593, N393, N607);
  and AND2_139 (keyinput_Wire_0[92], N354, N620);
  xor keyGate_0_92(N692, keyinput92, keyinput_Wire_0[92]);
  and AND2_140 (keyinput_Wire_0[93], N367, N620);
  xnor keyGate_0_93(KeyNOTWire_0[54], keyinput93, keyinput_Wire_0[93]);
  not KeyNOTGate_0_54(N693, KeyNOTWire_0[54]);
and AND2_141 (N694, N380, N620);
and AND2_142 (N695, N393, N620);
and AND2_143 (N696, N354, N625);
and AND2_144 (N697, N367, N625);
and AND2_145 (N698, N380, N625);
  and AND2_146 (keyinput_Wire_0[94], N393, N625);
  xor keyGate_0_94(KeyNOTWire_0[55], keyinput94, keyinput_Wire_0[94]);
  not KeyNOTGate_0_55(N699, KeyNOTWire_0[55]);
and AND2_147 (N700, N354, N630);
and AND2_148 (N701, N367, N630);
and AND2_149 (N702, N380, N630);
  and AND2_150 (keyinput_Wire_0[95], N393, N630);
  xor keyGate_0_95(N703, keyinput95, keyinput_Wire_0[95]);
  and AND2_151 (keyinput_Wire_0[96], N354, N635);
  xor keyGate_0_96(KeyNOTWire_0[56], keyinput96, keyinput_Wire_0[96]);
  not KeyNOTGate_0_56(N704, KeyNOTWire_0[56]);
and AND2_152 (N705, N367, N635);
  and AND2_153 (keyinput_Wire_0[97], N380, N635);
  xnor keyGate_0_97(N706, keyinput97, keyinput_Wire_0[97]);
and AND2_154 (N707, N393, N635);
  and AND2_155 (keyinput_Wire_0[98], N406, N640);
  xor keyGate_0_98(KeyNOTWire_0[57], keyinput98, keyinput_Wire_0[98]);
  not KeyNOTGate_0_57(N708, KeyNOTWire_0[57]);
  and AND2_156 (keyinput_Wire_0[99], N419, N640);
  xor keyGate_0_99(N709, keyinput99, keyinput_Wire_0[99]);
  and AND2_157 (keyinput_Wire_0[100], N432, N640);
  xor keyGate_0_100(N710, keyinput100, keyinput_Wire_0[100]);
and AND2_158 (N711, N445, N640);
  and AND2_159 (keyinput_Wire_0[101], N406, N645);
  xnor keyGate_0_101(KeyNOTWire_0[58], keyinput101, keyinput_Wire_0[101]);
  not KeyNOTGate_0_58(N712, KeyNOTWire_0[58]);
and AND2_160 (N713, N419, N645);
and AND2_161 (N714, N432, N645);
  and AND2_162 (keyinput_Wire_0[102], N445, N645);
  xor keyGate_0_102(N715, keyinput102, keyinput_Wire_0[102]);
  and AND2_163 (keyinput_Wire_0[103], N406, N650);
  xor keyGate_0_103(N716, keyinput103, keyinput_Wire_0[103]);
and AND2_164 (N717, N419, N650);
and AND2_165 (N718, N432, N650);
  and AND2_166 (keyinput_Wire_0[104], N445, N650);
  xor keyGate_0_104(N719, keyinput104, keyinput_Wire_0[104]);
and AND2_167 (N720, N406, N655);
  and AND2_168 (keyinput_Wire_0[105], N419, N655);
  xor keyGate_0_105(KeyNOTWire_0[59], keyinput105, keyinput_Wire_0[105]);
  not KeyNOTGate_0_59(N721, KeyNOTWire_0[59]);
  and AND2_169 (keyinput_Wire_0[106], N432, N655);
  xnor keyGate_0_106(KeyNOTWire_0[60], keyinput106, keyinput_Wire_0[106]);
  not KeyNOTGate_0_60(N722, KeyNOTWire_0[60]);
  and AND2_170 (keyinput_Wire_0[107], N445, N655);
  xor keyGate_0_107(N723, keyinput107, keyinput_Wire_0[107]);
  xor XOR2_171 (keyinput_Wire_0[108], N1, N692);
  xor keyGate_0_108(N724, keyinput108, keyinput_Wire_0[108]);
  xor XOR2_172 (keyinput_Wire_0[109], N5, N693);
  xnor keyGate_0_109(KeyNOTWire_0[61], keyinput109, keyinput_Wire_0[109]);
  not KeyNOTGate_0_61(N725, KeyNOTWire_0[61]);
  xor XOR2_173 (keyinput_Wire_0[110], N9, N694);
  xnor keyGate_0_110(KeyNOTWire_0[62], keyinput110, keyinput_Wire_0[110]);
  not KeyNOTGate_0_62(N726, KeyNOTWire_0[62]);
  xor XOR2_174 (keyinput_Wire_0[111], N13, N695);
  xor keyGate_0_111(N727, keyinput111, keyinput_Wire_0[111]);
  xor XOR2_175 (keyinput_Wire_0[112], N17, N696);
  xor keyGate_0_112(KeyNOTWire_0[63], keyinput112, keyinput_Wire_0[112]);
  not KeyNOTGate_0_63(N728, KeyNOTWire_0[63]);
  xor XOR2_176 (keyinput_Wire_0[113], N21, N697);
  xor keyGate_0_113(KeyNOTWire_0[64], keyinput113, keyinput_Wire_0[113]);
  not KeyNOTGate_0_64(N729, KeyNOTWire_0[64]);
xor XOR2_177 (N730, N25, N698);
xor XOR2_178 (N731, N29, N699);
  xor XOR2_179 (keyinput_Wire_0[114], N33, N700);
  xnor keyGate_0_114(N732, keyinput114, keyinput_Wire_0[114]);
  xor XOR2_180 (keyinput_Wire_0[115], N37, N701);
  xnor keyGate_0_115(KeyNOTWire_0[65], keyinput115, keyinput_Wire_0[115]);
  not KeyNOTGate_0_65(N733, KeyNOTWire_0[65]);
xor XOR2_181 (N734, N41, N702);
  xor XOR2_182 (keyinput_Wire_0[116], N45, N703);
  xnor keyGate_0_116(N735, keyinput116, keyinput_Wire_0[116]);
  xor XOR2_183 (keyinput_Wire_0[117], N49, N704);
  xnor keyGate_0_117(N736, keyinput117, keyinput_Wire_0[117]);
xor XOR2_184 (N737, N53, N705);
  xor XOR2_185 (keyinput_Wire_0[118], N57, N706);
  xnor keyGate_0_118(N738, keyinput118, keyinput_Wire_0[118]);
xor XOR2_186 (N739, N61, N707);
  xor XOR2_187 (keyinput_Wire_0[119], N65, N708);
  xor keyGate_0_119(N740, keyinput119, keyinput_Wire_0[119]);
  xor XOR2_188 (keyinput_Wire_0[120], N69, N709);
  xor keyGate_0_120(KeyNOTWire_0[66], keyinput120, keyinput_Wire_0[120]);
  not KeyNOTGate_0_66(N741, KeyNOTWire_0[66]);
  xor XOR2_189 (keyinput_Wire_0[121], N73, N710);
  xnor keyGate_0_121(KeyNOTWire_0[67], keyinput121, keyinput_Wire_0[121]);
  not KeyNOTGate_0_67(N742, KeyNOTWire_0[67]);
  xor XOR2_190 (keyinput_Wire_0[122], N77, N711);
  xnor keyGate_0_122(N743, keyinput122, keyinput_Wire_0[122]);
  xor XOR2_191 (keyinput_Wire_0[123], N81, N712);
  xnor keyGate_0_123(KeyNOTWire_0[68], keyinput123, keyinput_Wire_0[123]);
  not KeyNOTGate_0_68(N744, KeyNOTWire_0[68]);
  xor XOR2_192 (keyinput_Wire_0[124], N85, N713);
  xor keyGate_0_124(KeyNOTWire_0[69], keyinput124, keyinput_Wire_0[124]);
  not KeyNOTGate_0_69(N745, KeyNOTWire_0[69]);
xor XOR2_193 (N746, N89, N714);
xor XOR2_194 (N747, N93, N715);
xor XOR2_195 (N748, N97, N716);
  xor XOR2_196 (keyinput_Wire_0[125], N101, N717);
  xnor keyGate_0_125(N749, keyinput125, keyinput_Wire_0[125]);
  xor XOR2_197 (keyinput_Wire_0[126], N105, N718);
  xnor keyGate_0_126(KeyNOTWire_0[70], keyinput126, keyinput_Wire_0[126]);
  not KeyNOTGate_0_70(KeyWire_0_1, KeyNOTWire_0[70]);
  xor flip_it (N750, KeyWire_0_1, KeyWire_0_2 );
xor XOR2_198 (N751, N109, N719);
xor XOR2_199 (N752, N113, N720);
xor XOR2_200 (N753, N117, N721);
xor XOR2_201 (N754, N121, N722);
  xor XOR2_202 (keyinput_Wire_0[127], N125, N723);
  xor keyGate_0_127(N755, keyinput127, keyinput_Wire_0[127]);

AntiSAT some_name( KeyWire_0_2, N61, N137, N117, N129, N45, N125, N101, N37, N134, N105, N81, N136, N130, N29, N1, N41, N13, N53, N109, N69, N73, N85, N5, N131, N93, N49, N133, N89, N21, N33, N57, N113, N77, N65, N135, N25, N121, N132, N17, N97, N9, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
       keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
       keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
       keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
       keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
       keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
       keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
       keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
       keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
       keyinput250);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N61, N137, N117, N129, N45, N125, N101, N37, N134, N105, N81, N136, N130, N29, N1, N41, N13, N53, N109, N69, N73, N85, N5, N131, N93, N49, N133, N89, N21, N33, N57, N113, N77, N65, N135, N25, N121, N132, N17, N97, N9, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, keyinput208, keyinput209 ,
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
        keyinput250);

  input keyinput210, keyinput211, keyinput212, keyinput213, keyinput214;
  input keyinput215, keyinput216, keyinput217, keyinput218, keyinput219;
  input keyinput220, keyinput221, keyinput222, keyinput223, keyinput224;
  input keyinput225, keyinput226, keyinput227, keyinput228, keyinput229;
  input keyinput230, keyinput231, keyinput232, keyinput233, keyinput234;
  input keyinput235, keyinput236, keyinput237, keyinput238, keyinput239;
  input keyinput240, keyinput241, keyinput242, keyinput243, keyinput244;
  input keyinput245, keyinput246, keyinput247, keyinput248, keyinput249;
  input keyinput250;

  wire [0:40] keyNTin_Wire_1;
  wire [0:17] KeyNOTWire_1;

  input N61, N137, N117, N129, N45, N125, N101, N37, N134, N105, N81, N136, N130, N29, N1, N41, N13, N53, N109, N69, N73, N85, N5, N131, N93, N49, N133, N89, N21, N33, N57, N113, N77, N65, N135, N25, N121, N132, N17, N97, N9;
  input keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, keyinput208, keyinput209;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83 ;

  xnor KeyGate0 (newWire_0, N61, keyinput128);
  xnor KeyGate1 (newWire_1, N137, keyinput129);
  xnor KeyGate2 (newWire_2, N117, keyinput130);
  xor  KeyGate3 (keyNTin_Wire_1[0], N129, keyinput131);
  xor keyNTinGate_1_0(newWire_3, keyinput210, keyNTin_Wire_1[0]);
  xnor KeyGate4 (newWire_4, N45, keyinput132);
  xor  KeyGate5 (newWire_5, N125, keyinput133);
  xnor KeyGate6 (newWire_6, N101, keyinput134);
  xor  KeyGate7 (newWire_7, N37, keyinput135);
  xnor KeyGate8 (keyNTin_Wire_1[1], N134, keyinput136);
  xnor keyNTinGate_1_1(KeyNOTWire_1[0], keyinput211, keyNTin_Wire_1[1]);
  not KeyNOTGate_1_0(newWire_8, KeyNOTWire_1[0]);
  xnor KeyGate9 (newWire_9, N105, keyinput137);
  xnor KeyGate10 (keyNTin_Wire_1[2], N81, keyinput138);
  xnor keyNTinGate_1_2(KeyNOTWire_1[1], keyinput212, keyNTin_Wire_1[2]);
  not KeyNOTGate_1_1(newWire_10, KeyNOTWire_1[1]);
  xor  KeyGate11 (newWire_11, N136, keyinput139);
  xor  KeyGate12 (keyNTin_Wire_1[3], N130, keyinput140);
  xnor keyNTinGate_1_3(KeyNOTWire_1[2], keyinput213, keyNTin_Wire_1[3]);
  not KeyNOTGate_1_2(newWire_12, KeyNOTWire_1[2]);
  xor  KeyGate13 (keyNTin_Wire_1[4], N29, keyinput141);
  xor keyNTinGate_1_4(newWire_13, keyinput214, keyNTin_Wire_1[4]);
  xnor KeyGate14 (newWire_14, N1, keyinput142);
  xnor KeyGate15 (newWire_15, N41, keyinput143);
  xnor KeyGate16 (keyNTin_Wire_1[5], N13, keyinput144);
  xor keyNTinGate_1_5(KeyNOTWire_1[3], keyinput215, keyNTin_Wire_1[5]);
  not KeyNOTGate_1_3(newWire_16, KeyNOTWire_1[3]);
  xor  KeyGate17 (newWire_17, N53, keyinput145);
  xor  KeyGate18 (keyNTin_Wire_1[6], N109, keyinput146);
  xnor keyNTinGate_1_6(KeyNOTWire_1[4], keyinput216, keyNTin_Wire_1[6]);
  not KeyNOTGate_1_4(newWire_18, KeyNOTWire_1[4]);
  xnor KeyGate19 (keyNTin_Wire_1[7], N69, keyinput147);
  xnor keyNTinGate_1_7(KeyNOTWire_1[5], keyinput217, keyNTin_Wire_1[7]);
  not KeyNOTGate_1_5(newWire_19, KeyNOTWire_1[5]);
  xor  KeyGate20 (keyNTin_Wire_1[8], N73, keyinput148);
  xnor keyNTinGate_1_8(newWire_20, keyinput218, keyNTin_Wire_1[8]);
  xor  KeyGate21 (newWire_21, N85, keyinput149);
  xor  KeyGate22 (newWire_22, N5, keyinput150);
  xor  KeyGate23 (keyNTin_Wire_1[9], N131, keyinput151);
  xnor keyNTinGate_1_9(KeyNOTWire_1[6], keyinput219, keyNTin_Wire_1[9]);
  not KeyNOTGate_1_6(newWire_23, KeyNOTWire_1[6]);
  xnor KeyGate24 (newWire_24, N93, keyinput152);
  xor  KeyGate25 (keyNTin_Wire_1[10], N49, keyinput153);
  xor keyNTinGate_1_10(KeyNOTWire_1[7], keyinput220, keyNTin_Wire_1[10]);
  not KeyNOTGate_1_7(newWire_25, KeyNOTWire_1[7]);
  xnor KeyGate26 (newWire_26, N133, keyinput154);
  xnor KeyGate27 (newWire_27, N89, keyinput155);
  xor  KeyGate28 (keyNTin_Wire_1[11], N21, keyinput156);
  xnor keyNTinGate_1_11(newWire_28, keyinput221, keyNTin_Wire_1[11]);
  xor  KeyGate29 (keyNTin_Wire_1[12], N33, keyinput157);
  xnor keyNTinGate_1_12(KeyNOTWire_1[8], keyinput222, keyNTin_Wire_1[12]);
  not KeyNOTGate_1_8(newWire_29, KeyNOTWire_1[8]);
  xnor KeyGate30 (newWire_30, N57, keyinput158);
  xor  KeyGate31 (newWire_31, N113, keyinput159);
  xnor KeyGate32 (newWire_32, N77, keyinput160);
  xor  KeyGate33 (newWire_33, N65, keyinput161);
  xor  KeyGate34 (keyNTin_Wire_1[13], N135, keyinput162);
  xnor keyNTinGate_1_13(KeyNOTWire_1[9], keyinput223, keyNTin_Wire_1[13]);
  not KeyNOTGate_1_9(newWire_34, KeyNOTWire_1[9]);
  xor  KeyGate35 (newWire_35, N25, keyinput163);
  xor  KeyGate36 (keyNTin_Wire_1[14], N121, keyinput164);
  xor keyNTinGate_1_14(KeyNOTWire_1[10], keyinput224, keyNTin_Wire_1[14]);
  not KeyNOTGate_1_10(newWire_36, KeyNOTWire_1[10]);
  xnor KeyGate37 (keyNTin_Wire_1[15], N132, keyinput165);
  xor keyNTinGate_1_15(KeyNOTWire_1[11], keyinput225, keyNTin_Wire_1[15]);
  not KeyNOTGate_1_11(newWire_37, KeyNOTWire_1[11]);
  xor  KeyGate38 (newWire_38, N17, keyinput166);
  xnor KeyGate39 (newWire_39, N97, keyinput167);
  xnor KeyGate40 (keyNTin_Wire_1[16], N9, keyinput168);
  xnor keyNTinGate_1_16(newWire_40, keyinput226, keyNTin_Wire_1[16]);
  xnor KeyGate41 (newWire_41, N61, keyinput169);
  xnor KeyGate42 (newWire_42, N137, keyinput170);
  xnor KeyGate43 (keyNTin_Wire_1[17], N117, keyinput171);
  xor keyNTinGate_1_17(KeyNOTWire_1[12], keyinput227, keyNTin_Wire_1[17]);
  not KeyNOTGate_1_12(newWire_43, KeyNOTWire_1[12]);
  xor  KeyGate44 (keyNTin_Wire_1[18], N129, keyinput172);
  xor keyNTinGate_1_18(KeyNOTWire_1[13], keyinput228, keyNTin_Wire_1[18]);
  not KeyNOTGate_1_13(newWire_44, KeyNOTWire_1[13]);
  xnor KeyGate45 (keyNTin_Wire_1[19], N45, keyinput173);
  xnor keyNTinGate_1_19(newWire_45, keyinput229, keyNTin_Wire_1[19]);
  xnor KeyGate46 (newWire_46, N125, keyinput174);
  xnor KeyGate47 (newWire_47, N101, keyinput175);
  xor  KeyGate48 (newWire_48, N37, keyinput176);
  xnor KeyGate49 (newWire_49, N134, keyinput177);
  xor  KeyGate50 (keyNTin_Wire_1[20], N105, keyinput178);
  xnor keyNTinGate_1_20(KeyNOTWire_1[14], keyinput230, keyNTin_Wire_1[20]);
  not KeyNOTGate_1_14(newWire_50, KeyNOTWire_1[14]);
  xor  KeyGate51 (keyNTin_Wire_1[21], N81, keyinput179);
  xor keyNTinGate_1_21(newWire_51, keyinput231, keyNTin_Wire_1[21]);
  xnor KeyGate52 (newWire_52, N136, keyinput180);
  xnor KeyGate53 (keyNTin_Wire_1[22], N130, keyinput181);
  xor keyNTinGate_1_22(newWire_53, keyinput232, keyNTin_Wire_1[22]);
  xor  KeyGate54 (newWire_54, N29, keyinput182);
  xnor KeyGate55 (keyNTin_Wire_1[23], N1, keyinput183);
  xor keyNTinGate_1_23(newWire_55, keyinput233, keyNTin_Wire_1[23]);
  xor  KeyGate56 (keyNTin_Wire_1[24], N41, keyinput184);
  xnor keyNTinGate_1_24(newWire_56, keyinput234, keyNTin_Wire_1[24]);
  xor  KeyGate57 (newWire_57, N13, keyinput185);
  xnor KeyGate58 (keyNTin_Wire_1[25], N53, keyinput186);
  xnor keyNTinGate_1_25(KeyNOTWire_1[15], keyinput235, keyNTin_Wire_1[25]);
  not KeyNOTGate_1_15(newWire_58, KeyNOTWire_1[15]);
  xor  KeyGate59 (keyNTin_Wire_1[26], N109, keyinput187);
  xor keyNTinGate_1_26(newWire_59, keyinput236, keyNTin_Wire_1[26]);
  xor  KeyGate60 (keyNTin_Wire_1[27], N69, keyinput188);
  xnor keyNTinGate_1_27(KeyNOTWire_1[16], keyinput237, keyNTin_Wire_1[27]);
  not KeyNOTGate_1_16(newWire_60, KeyNOTWire_1[16]);
  xnor KeyGate61 (keyNTin_Wire_1[28], N73, keyinput189);
  xnor keyNTinGate_1_28(newWire_61, keyinput238, keyNTin_Wire_1[28]);
  xnor KeyGate62 (keyNTin_Wire_1[29], N85, keyinput190);
  xor keyNTinGate_1_29(newWire_62, keyinput239, keyNTin_Wire_1[29]);
  xor  KeyGate63 (newWire_63, N5, keyinput191);
  xnor KeyGate64 (keyNTin_Wire_1[30], N131, keyinput192);
  xor keyNTinGate_1_30(newWire_64, keyinput240, keyNTin_Wire_1[30]);
  xnor KeyGate65 (newWire_65, N93, keyinput193);
  xnor KeyGate66 (keyNTin_Wire_1[31], N49, keyinput194);
  xnor keyNTinGate_1_31(newWire_66, keyinput241, keyNTin_Wire_1[31]);
  xor  KeyGate67 (newWire_67, N133, keyinput195);
  xnor KeyGate68 (newWire_68, N89, keyinput196);
  xnor KeyGate69 (newWire_69, N21, keyinput197);
  xnor KeyGate70 (keyNTin_Wire_1[32], N33, keyinput198);
  xnor keyNTinGate_1_32(newWire_70, keyinput242, keyNTin_Wire_1[32]);
  xor  KeyGate71 (newWire_71, N57, keyinput199);
  xnor KeyGate72 (keyNTin_Wire_1[33], N113, keyinput200);
  xnor keyNTinGate_1_33(newWire_72, keyinput243, keyNTin_Wire_1[33]);
  xor  KeyGate73 (keyNTin_Wire_1[34], N77, keyinput201);
  xnor keyNTinGate_1_34(newWire_73, keyinput244, keyNTin_Wire_1[34]);
  xor  KeyGate74 (newWire_74, N65, keyinput202);
  xnor KeyGate75 (newWire_75, N135, keyinput203);
  xor  KeyGate76 (keyNTin_Wire_1[35], N25, keyinput204);
  xor keyNTinGate_1_35(newWire_76, keyinput245, keyNTin_Wire_1[35]);
  xnor KeyGate77 (keyNTin_Wire_1[36], N121, keyinput205);
  xor keyNTinGate_1_36(newWire_77, keyinput246, keyNTin_Wire_1[36]);
  xnor KeyGate78 (newWire_78, N132, keyinput206);
  xor  KeyGate79 (keyNTin_Wire_1[37], N17, keyinput207);
  xnor keyNTinGate_1_37(KeyNOTWire_1[17], keyinput247, keyNTin_Wire_1[37]);
  not KeyNOTGate_1_17(newWire_79, KeyNOTWire_1[17]);
  xor  KeyGate80 (keyNTin_Wire_1[38], N97, keyinput208);
  xor keyNTinGate_1_38(newWire_80, keyinput248, keyNTin_Wire_1[38]);
  xor  KeyGate81 (newWire_81, N9, keyinput209);
  and some_function (keyNTin_Wire_1[39], newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40 );
  xor keyNTinGate_1_39(newWire_82, keyinput249, keyNTin_Wire_1[39]);
  nand compl_function (newWire_83, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81);
  and finalAND (keyNTin_Wire_1[40], newWire_82, newWire_83);
  xnor keyNTinGate_1_40(KeyWire_0_2, keyinput250, keyNTin_Wire_1[40]);

endmodule /* AntiSAT */
