`timescale 1ns / 1ps
// Verilog
// c432
// Ninputs 36
// Noutputs 7
// NtotalGates 160
// NOT1 40
// NAND2 64
// NOR2 19
// AND9 3
// XOR2 18
// NAND4 14
// AND8 1
// NAND3 1

module top (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
                  N430,N431,N432,
        keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4,
        keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9,
        keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14,
        keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19,
        keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24,
        keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29,
        keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34,
        keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39,
        keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44,
        keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49,
        keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54,
        keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59,
        keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64,
        keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69,
        keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74,
        keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79,
        keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84,
        keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89,
        keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94,
        keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99,
        keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104,
        keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109,
        keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114,
        keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119,
        keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124,
        keyIn_0_125, keyIn_0_126, keyIn_0_127);

  input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4;
  input keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9;
  input keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14;
  input keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19;
  input keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24;
  input keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29;
  input keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34;
  input keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39;
  input keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44;
  input keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49;
  input keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54;
  input keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59;
  input keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64;
  input keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69;
  input keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74;
  input keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79;
  input keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84;
  input keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89;
  input keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94;
  input keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99;
  input keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104;
  input keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109;
  input keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114;
  input keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119;
  input keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124;
  input keyIn_0_125, keyIn_0_126, keyIn_0_127;

  wire [0:127] KeyWire_0;
  wire [0:56] KeyNOTWire_0;

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;

output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429;

  not NOT1_1 (KeyWire_0[0], N1);
  xnor KeyGate_0_0(N118, keyIn_0_0, KeyWire_0[0]);
  not NOT1_2 (KeyWire_0[1], N4);
  xnor KeyGate_0_1(N119, keyIn_0_1, KeyWire_0[1]);
  not NOT1_3 (KeyWire_0[2], N11);
  xor KeyGate_0_2(N122, keyIn_0_2, KeyWire_0[2]);
  not NOT1_4 (KeyWire_0[3], N17);
  xor KeyGate_0_3(KeyNOTWire_0[0], keyIn_0_3, KeyWire_0[3]);
  not KeyNOTGate_0_0(N123, KeyNOTWire_0[0]);
  not NOT1_5 (KeyWire_0[4], N24);
  xor KeyGate_0_4(N126, keyIn_0_4, KeyWire_0[4]);
  not NOT1_6 (KeyWire_0[5], N30);
  xor KeyGate_0_5(KeyNOTWire_0[1], keyIn_0_5, KeyWire_0[5]);
  not KeyNOTGate_0_1(N127, KeyNOTWire_0[1]);
  not NOT1_7 (KeyWire_0[6], N37);
  xnor KeyGate_0_6(KeyNOTWire_0[2], keyIn_0_6, KeyWire_0[6]);
  not KeyNOTGate_0_2(N130, KeyNOTWire_0[2]);
  not NOT1_8 (KeyWire_0[7], N43);
  xnor KeyGate_0_7(KeyNOTWire_0[3], keyIn_0_7, KeyWire_0[7]);
  not KeyNOTGate_0_3(N131, KeyNOTWire_0[3]);
  not NOT1_9 (KeyWire_0[8], N50);
  xor KeyGate_0_8(N134, keyIn_0_8, KeyWire_0[8]);
  not NOT1_10 (KeyWire_0[9], N56);
  xor KeyGate_0_9(N135, keyIn_0_9, KeyWire_0[9]);
  not NOT1_11 (KeyWire_0[10], N63);
  xor KeyGate_0_10(KeyNOTWire_0[4], keyIn_0_10, KeyWire_0[10]);
  not KeyNOTGate_0_4(N138, KeyNOTWire_0[4]);
  not NOT1_12 (KeyWire_0[11], N69);
  xnor KeyGate_0_11(KeyNOTWire_0[5], keyIn_0_11, KeyWire_0[11]);
  not KeyNOTGate_0_5(N139, KeyNOTWire_0[5]);
  not NOT1_13 (KeyWire_0[12], N76);
  xnor KeyGate_0_12(N142, keyIn_0_12, KeyWire_0[12]);
  not NOT1_14 (KeyWire_0[13], N82);
  xnor KeyGate_0_13(N143, keyIn_0_13, KeyWire_0[13]);
  not NOT1_15 (KeyWire_0[14], N89);
  xnor KeyGate_0_14(KeyNOTWire_0[6], keyIn_0_14, KeyWire_0[14]);
  not KeyNOTGate_0_6(N146, KeyNOTWire_0[6]);
  not NOT1_16 (KeyWire_0[15], N95);
  xnor KeyGate_0_15(KeyNOTWire_0[7], keyIn_0_15, KeyWire_0[15]);
  not KeyNOTGate_0_7(N147, KeyNOTWire_0[7]);
  not NOT1_17 (KeyWire_0[16], N102);
  xor KeyGate_0_16(N150, keyIn_0_16, KeyWire_0[16]);
  not NOT1_18 (KeyWire_0[17], N108);
  xnor KeyGate_0_17(N151, keyIn_0_17, KeyWire_0[17]);
  nand NAND2_19 (KeyWire_0[18], N118, N4);
  xnor KeyGate_0_18(KeyNOTWire_0[8], keyIn_0_18, KeyWire_0[18]);
  not KeyNOTGate_0_8(N154, KeyNOTWire_0[8]);
  nor NOR2_20 (KeyWire_0[19], N8, N119);
  xnor KeyGate_0_19(KeyNOTWire_0[9], keyIn_0_19, KeyWire_0[19]);
  not KeyNOTGate_0_9(N157, KeyNOTWire_0[9]);
nor NOR2_21 (N158, N14, N119);
  nand NAND2_22 (KeyWire_0[20], N122, N17);
  xor KeyGate_0_20(N159, keyIn_0_20, KeyWire_0[20]);
  nand NAND2_23 (KeyWire_0[21], N126, N30);
  xor KeyGate_0_21(KeyNOTWire_0[10], keyIn_0_21, KeyWire_0[21]);
  not KeyNOTGate_0_10(N162, KeyNOTWire_0[10]);
  nand NAND2_24 (KeyWire_0[22], N130, N43);
  xor KeyGate_0_22(N165, keyIn_0_22, KeyWire_0[22]);
  nand NAND2_25 (KeyWire_0[23], N134, N56);
  xor KeyGate_0_23(KeyNOTWire_0[11], keyIn_0_23, KeyWire_0[23]);
  not KeyNOTGate_0_11(N168, KeyNOTWire_0[11]);
  nand NAND2_26 (KeyWire_0[24], N138, N69);
  xnor KeyGate_0_24(N171, keyIn_0_24, KeyWire_0[24]);
  nand NAND2_27 (KeyWire_0[25], N142, N82);
  xor KeyGate_0_25(N174, keyIn_0_25, KeyWire_0[25]);
  nand NAND2_28 (KeyWire_0[26], N146, N95);
  xnor KeyGate_0_26(N177, keyIn_0_26, KeyWire_0[26]);
  nand NAND2_29 (KeyWire_0[27], N150, N108);
  xor KeyGate_0_27(N180, keyIn_0_27, KeyWire_0[27]);
  nor NOR2_30 (KeyWire_0[28], N21, N123);
  xor KeyGate_0_28(KeyNOTWire_0[12], keyIn_0_28, KeyWire_0[28]);
  not KeyNOTGate_0_12(N183, KeyNOTWire_0[12]);
nor NOR2_31 (N184, N27, N123);
  nor NOR2_32 (KeyWire_0[29], N34, N127);
  xor KeyGate_0_29(KeyNOTWire_0[13], keyIn_0_29, KeyWire_0[29]);
  not KeyNOTGate_0_13(N185, KeyNOTWire_0[13]);
nor NOR2_33 (N186, N40, N127);
  nor NOR2_34 (KeyWire_0[30], N47, N131);
  xor KeyGate_0_30(KeyNOTWire_0[14], keyIn_0_30, KeyWire_0[30]);
  not KeyNOTGate_0_14(N187, KeyNOTWire_0[14]);
nor NOR2_35 (N188, N53, N131);
  nor NOR2_36 (KeyWire_0[31], N60, N135);
  xnor KeyGate_0_31(N189, keyIn_0_31, KeyWire_0[31]);
nor NOR2_37 (N190, N66, N135);
  nor NOR2_38 (KeyWire_0[32], N73, N139);
  xor KeyGate_0_32(N191, keyIn_0_32, KeyWire_0[32]);
nor NOR2_39 (N192, N79, N139);
  nor NOR2_40 (KeyWire_0[33], N86, N143);
  xnor KeyGate_0_33(KeyNOTWire_0[15], keyIn_0_33, KeyWire_0[33]);
  not KeyNOTGate_0_15(N193, KeyNOTWire_0[15]);
nor NOR2_41 (N194, N92, N143);
  nor NOR2_42 (KeyWire_0[34], N99, N147);
  xor KeyGate_0_34(N195, keyIn_0_34, KeyWire_0[34]);
nor NOR2_43 (N196, N105, N147);
  nor NOR2_44 (KeyWire_0[35], N112, N151);
  xor KeyGate_0_35(KeyNOTWire_0[16], keyIn_0_35, KeyWire_0[35]);
  not KeyNOTGate_0_16(N197, KeyNOTWire_0[16]);
nor NOR2_45 (N198, N115, N151);
  and AND9_46 (KeyWire_0[36], N154, N159, N162, N165, N168, N171, N174, N177, N180);
  xnor KeyGate_0_36(KeyNOTWire_0[17], keyIn_0_36, KeyWire_0[36]);
  not KeyNOTGate_0_17(N199, KeyNOTWire_0[17]);
  not NOT1_47 (KeyWire_0[37], N199);
  xnor KeyGate_0_37(KeyNOTWire_0[18], keyIn_0_37, KeyWire_0[37]);
  not KeyNOTGate_0_18(N203, KeyNOTWire_0[18]);
not NOT1_48 (N213, N199);
not NOT1_49 (N223, N199);
  xor XOR2_50 (KeyWire_0[38], N203, N154);
  xor KeyGate_0_38(KeyNOTWire_0[19], keyIn_0_38, KeyWire_0[38]);
  not KeyNOTGate_0_19(N224, KeyNOTWire_0[19]);
  xor XOR2_51 (KeyWire_0[39], N203, N159);
  xor KeyGate_0_39(KeyNOTWire_0[20], keyIn_0_39, KeyWire_0[39]);
  not KeyNOTGate_0_20(N227, KeyNOTWire_0[20]);
  xor XOR2_52 (KeyWire_0[40], N203, N162);
  xnor KeyGate_0_40(N230, keyIn_0_40, KeyWire_0[40]);
  xor XOR2_53 (KeyWire_0[41], N203, N165);
  xor KeyGate_0_41(N233, keyIn_0_41, KeyWire_0[41]);
  xor XOR2_54 (KeyWire_0[42], N203, N168);
  xor KeyGate_0_42(N236, keyIn_0_42, KeyWire_0[42]);
  xor XOR2_55 (KeyWire_0[43], N203, N171);
  xnor KeyGate_0_43(N239, keyIn_0_43, KeyWire_0[43]);
nand NAND2_56 (N242, N1, N213);
  xor XOR2_57 (KeyWire_0[44], N203, N174);
  xor KeyGate_0_44(N243, keyIn_0_44, KeyWire_0[44]);
  nand NAND2_58 (KeyWire_0[45], N213, N11);
  xor KeyGate_0_45(KeyNOTWire_0[21], keyIn_0_45, KeyWire_0[45]);
  not KeyNOTGate_0_21(N246, KeyNOTWire_0[21]);
  xor XOR2_59 (KeyWire_0[46], N203, N177);
  xor KeyGate_0_46(N247, keyIn_0_46, KeyWire_0[46]);
nand NAND2_60 (N250, N213, N24);
  xor XOR2_61 (KeyWire_0[47], N203, N180);
  xnor KeyGate_0_47(KeyNOTWire_0[22], keyIn_0_47, KeyWire_0[47]);
  not KeyNOTGate_0_22(N251, KeyNOTWire_0[22]);
nand NAND2_62 (N254, N213, N37);
nand NAND2_63 (N255, N213, N50);
nand NAND2_64 (N256, N213, N63);
nand NAND2_65 (N257, N213, N76);
nand NAND2_66 (N258, N213, N89);
nand NAND2_67 (N259, N213, N102);
  nand NAND2_68 (KeyWire_0[48], N224, N157);
  xnor KeyGate_0_48(N260, keyIn_0_48, KeyWire_0[48]);
nand NAND2_69 (N263, N224, N158);
  nand NAND2_70 (KeyWire_0[49], N227, N183);
  xor KeyGate_0_49(N264, keyIn_0_49, KeyWire_0[49]);
  nand NAND2_71 (KeyWire_0[50], N230, N185);
  xnor KeyGate_0_50(N267, keyIn_0_50, KeyWire_0[50]);
  nand NAND2_72 (KeyWire_0[51], N233, N187);
  xnor KeyGate_0_51(KeyNOTWire_0[23], keyIn_0_51, KeyWire_0[51]);
  not KeyNOTGate_0_23(N270, KeyNOTWire_0[23]);
  nand NAND2_73 (KeyWire_0[52], N236, N189);
  xor KeyGate_0_52(KeyNOTWire_0[24], keyIn_0_52, KeyWire_0[52]);
  not KeyNOTGate_0_24(N273, KeyNOTWire_0[24]);
  nand NAND2_74 (KeyWire_0[53], N239, N191);
  xor KeyGate_0_53(N276, keyIn_0_53, KeyWire_0[53]);
  nand NAND2_75 (KeyWire_0[54], N243, N193);
  xnor KeyGate_0_54(N279, keyIn_0_54, KeyWire_0[54]);
  nand NAND2_76 (KeyWire_0[55], N247, N195);
  xor KeyGate_0_55(KeyNOTWire_0[25], keyIn_0_55, KeyWire_0[55]);
  not KeyNOTGate_0_25(N282, KeyNOTWire_0[25]);
  nand NAND2_77 (KeyWire_0[56], N251, N197);
  xnor KeyGate_0_56(N285, keyIn_0_56, KeyWire_0[56]);
nand NAND2_78 (N288, N227, N184);
nand NAND2_79 (N289, N230, N186);
nand NAND2_80 (N290, N233, N188);
  nand NAND2_81 (KeyWire_0[57], N236, N190);
  xnor KeyGate_0_57(N291, keyIn_0_57, KeyWire_0[57]);
  nand NAND2_82 (KeyWire_0[58], N239, N192);
  xnor KeyGate_0_58(KeyNOTWire_0[26], keyIn_0_58, KeyWire_0[58]);
  not KeyNOTGate_0_26(N292, KeyNOTWire_0[26]);
nand NAND2_83 (N293, N243, N194);
  nand NAND2_84 (KeyWire_0[59], N247, N196);
  xor KeyGate_0_59(N294, keyIn_0_59, KeyWire_0[59]);
nand NAND2_85 (N295, N251, N198);
  and AND9_86 (KeyWire_0[60], N260, N264, N267, N270, N273, N276, N279, N282, N285);
  xnor KeyGate_0_60(KeyNOTWire_0[27], keyIn_0_60, KeyWire_0[60]);
  not KeyNOTGate_0_27(N296, KeyNOTWire_0[27]);
not NOT1_87 (N300, N263);
not NOT1_88 (N301, N288);
not NOT1_89 (N302, N289);
not NOT1_90 (N303, N290);
  not NOT1_91 (KeyWire_0[61], N291);
  xnor KeyGate_0_61(N304, keyIn_0_61, KeyWire_0[61]);
  not NOT1_92 (KeyWire_0[62], N292);
  xnor KeyGate_0_62(N305, keyIn_0_62, KeyWire_0[62]);
not NOT1_93 (N306, N293);
  not NOT1_94 (KeyWire_0[63], N294);
  xor KeyGate_0_63(N307, keyIn_0_63, KeyWire_0[63]);
not NOT1_95 (N308, N295);
  not NOT1_96 (KeyWire_0[64], N296);
  xor KeyGate_0_64(N309, keyIn_0_64, KeyWire_0[64]);
  not NOT1_97 (KeyWire_0[65], N296);
  xor KeyGate_0_65(KeyNOTWire_0[28], keyIn_0_65, KeyWire_0[65]);
  not KeyNOTGate_0_28(N319, KeyNOTWire_0[28]);
not NOT1_98 (N329, N296);
  xor XOR2_99 (KeyWire_0[66], N309, N260);
  xor KeyGate_0_66(N330, keyIn_0_66, KeyWire_0[66]);
  xor XOR2_100 (KeyWire_0[67], N309, N264);
  xnor KeyGate_0_67(KeyNOTWire_0[29], keyIn_0_67, KeyWire_0[67]);
  not KeyNOTGate_0_29(N331, KeyNOTWire_0[29]);
  xor XOR2_101 (KeyWire_0[68], N309, N267);
  xnor KeyGate_0_68(N332, keyIn_0_68, KeyWire_0[68]);
  xor XOR2_102 (KeyWire_0[69], N309, N270);
  xnor KeyGate_0_69(KeyNOTWire_0[30], keyIn_0_69, KeyWire_0[69]);
  not KeyNOTGate_0_30(N333, KeyNOTWire_0[30]);
  nand NAND2_103 (KeyWire_0[70], N8, N319);
  xor KeyGate_0_70(N334, keyIn_0_70, KeyWire_0[70]);
  xor XOR2_104 (KeyWire_0[71], N309, N273);
  xnor KeyGate_0_71(KeyNOTWire_0[31], keyIn_0_71, KeyWire_0[71]);
  not KeyNOTGate_0_31(N335, KeyNOTWire_0[31]);
  nand NAND2_105 (KeyWire_0[72], N319, N21);
  xnor KeyGate_0_72(KeyNOTWire_0[32], keyIn_0_72, KeyWire_0[72]);
  not KeyNOTGate_0_32(N336, KeyNOTWire_0[32]);
  xor XOR2_106 (KeyWire_0[73], N309, N276);
  xor KeyGate_0_73(N337, keyIn_0_73, KeyWire_0[73]);
  nand NAND2_107 (KeyWire_0[74], N319, N34);
  xor KeyGate_0_74(N338, keyIn_0_74, KeyWire_0[74]);
  xor XOR2_108 (KeyWire_0[75], N309, N279);
  xor KeyGate_0_75(KeyNOTWire_0[33], keyIn_0_75, KeyWire_0[75]);
  not KeyNOTGate_0_33(N339, KeyNOTWire_0[33]);
  nand NAND2_109 (KeyWire_0[76], N319, N47);
  xor KeyGate_0_76(N340, keyIn_0_76, KeyWire_0[76]);
  xor XOR2_110 (KeyWire_0[77], N309, N282);
  xor KeyGate_0_77(N341, keyIn_0_77, KeyWire_0[77]);
  nand NAND2_111 (KeyWire_0[78], N319, N60);
  xnor KeyGate_0_78(N342, keyIn_0_78, KeyWire_0[78]);
  xor XOR2_112 (KeyWire_0[79], N309, N285);
  xnor KeyGate_0_79(N343, keyIn_0_79, KeyWire_0[79]);
  nand NAND2_113 (KeyWire_0[80], N319, N73);
  xnor KeyGate_0_80(KeyNOTWire_0[34], keyIn_0_80, KeyWire_0[80]);
  not KeyNOTGate_0_34(N344, KeyNOTWire_0[34]);
  nand NAND2_114 (KeyWire_0[81], N319, N86);
  xor KeyGate_0_81(N345, keyIn_0_81, KeyWire_0[81]);
  nand NAND2_115 (KeyWire_0[82], N319, N99);
  xnor KeyGate_0_82(N346, keyIn_0_82, KeyWire_0[82]);
  nand NAND2_116 (KeyWire_0[83], N319, N112);
  xor KeyGate_0_83(N347, keyIn_0_83, KeyWire_0[83]);
  nand NAND2_117 (KeyWire_0[84], N330, N300);
  xnor KeyGate_0_84(N348, keyIn_0_84, KeyWire_0[84]);
  nand NAND2_118 (KeyWire_0[85], N331, N301);
  xor KeyGate_0_85(N349, keyIn_0_85, KeyWire_0[85]);
  nand NAND2_119 (KeyWire_0[86], N332, N302);
  xnor KeyGate_0_86(KeyNOTWire_0[35], keyIn_0_86, KeyWire_0[86]);
  not KeyNOTGate_0_35(N350, KeyNOTWire_0[35]);
  nand NAND2_120 (KeyWire_0[87], N333, N303);
  xor KeyGate_0_87(KeyNOTWire_0[36], keyIn_0_87, KeyWire_0[87]);
  not KeyNOTGate_0_36(N351, KeyNOTWire_0[36]);
  nand NAND2_121 (KeyWire_0[88], N335, N304);
  xnor KeyGate_0_88(KeyNOTWire_0[37], keyIn_0_88, KeyWire_0[88]);
  not KeyNOTGate_0_37(N352, KeyNOTWire_0[37]);
  nand NAND2_122 (KeyWire_0[89], N337, N305);
  xor KeyGate_0_89(KeyNOTWire_0[38], keyIn_0_89, KeyWire_0[89]);
  not KeyNOTGate_0_38(N353, KeyNOTWire_0[38]);
  nand NAND2_123 (KeyWire_0[90], N339, N306);
  xor KeyGate_0_90(KeyNOTWire_0[39], keyIn_0_90, KeyWire_0[90]);
  not KeyNOTGate_0_39(N354, KeyNOTWire_0[39]);
  nand NAND2_124 (KeyWire_0[91], N341, N307);
  xor KeyGate_0_91(N355, keyIn_0_91, KeyWire_0[91]);
  nand NAND2_125 (KeyWire_0[92], N343, N308);
  xor KeyGate_0_92(KeyNOTWire_0[40], keyIn_0_92, KeyWire_0[92]);
  not KeyNOTGate_0_40(N356, KeyNOTWire_0[40]);
  and AND9_126 (KeyWire_0[93], N348, N349, N350, N351, N352, N353, N354, N355, N356);
  xor KeyGate_0_93(N357, keyIn_0_93, KeyWire_0[93]);
  not NOT1_127 (KeyWire_0[94], N357);
  xnor KeyGate_0_94(KeyNOTWire_0[41], keyIn_0_94, KeyWire_0[94]);
  not KeyNOTGate_0_41(N360, KeyNOTWire_0[41]);
  not NOT1_128 (KeyWire_0[95], N357);
  xnor KeyGate_0_95(KeyNOTWire_0[42], keyIn_0_95, KeyWire_0[95]);
  not KeyNOTGate_0_42(N370, KeyNOTWire_0[42]);
  nand NAND2_129 (KeyWire_0[96], N14, N360);
  xnor KeyGate_0_96(N371, keyIn_0_96, KeyWire_0[96]);
  nand NAND2_130 (KeyWire_0[97], N360, N27);
  xor KeyGate_0_97(KeyNOTWire_0[43], keyIn_0_97, KeyWire_0[97]);
  not KeyNOTGate_0_43(N372, KeyNOTWire_0[43]);
  nand NAND2_131 (KeyWire_0[98], N360, N40);
  xnor KeyGate_0_98(N373, keyIn_0_98, KeyWire_0[98]);
  nand NAND2_132 (KeyWire_0[99], N360, N53);
  xnor KeyGate_0_99(N374, keyIn_0_99, KeyWire_0[99]);
  nand NAND2_133 (KeyWire_0[100], N360, N66);
  xor KeyGate_0_100(N375, keyIn_0_100, KeyWire_0[100]);
  nand NAND2_134 (KeyWire_0[101], N360, N79);
  xor KeyGate_0_101(KeyNOTWire_0[44], keyIn_0_101, KeyWire_0[101]);
  not KeyNOTGate_0_44(N376, KeyNOTWire_0[44]);
  nand NAND2_135 (KeyWire_0[102], N360, N92);
  xor KeyGate_0_102(N377, keyIn_0_102, KeyWire_0[102]);
  nand NAND2_136 (KeyWire_0[103], N360, N105);
  xor KeyGate_0_103(KeyNOTWire_0[45], keyIn_0_103, KeyWire_0[103]);
  not KeyNOTGate_0_45(N378, KeyNOTWire_0[45]);
  nand NAND2_137 (KeyWire_0[104], N360, N115);
  xnor KeyGate_0_104(N379, keyIn_0_104, KeyWire_0[104]);
  nand NAND4_138 (KeyWire_0[105], N4, N242, N334, N371);
  xnor KeyGate_0_105(N380, keyIn_0_105, KeyWire_0[105]);
  nand NAND4_139 (KeyWire_0[106], N246, N336, N372, N17);
  xnor KeyGate_0_106(N381, keyIn_0_106, KeyWire_0[106]);
  nand NAND4_140 (KeyWire_0[107], N250, N338, N373, N30);
  xor KeyGate_0_107(KeyNOTWire_0[46], keyIn_0_107, KeyWire_0[107]);
  not KeyNOTGate_0_46(N386, KeyNOTWire_0[46]);
  nand NAND4_141 (KeyWire_0[108], N254, N340, N374, N43);
  xor KeyGate_0_108(N393, keyIn_0_108, KeyWire_0[108]);
  nand NAND4_142 (KeyWire_0[109], N255, N342, N375, N56);
  xnor KeyGate_0_109(N399, keyIn_0_109, KeyWire_0[109]);
  nand NAND4_143 (KeyWire_0[110], N256, N344, N376, N69);
  xor KeyGate_0_110(KeyNOTWire_0[47], keyIn_0_110, KeyWire_0[110]);
  not KeyNOTGate_0_47(N404, KeyNOTWire_0[47]);
  nand NAND4_144 (KeyWire_0[111], N257, N345, N377, N82);
  xor KeyGate_0_111(N407, keyIn_0_111, KeyWire_0[111]);
  nand NAND4_145 (KeyWire_0[112], N258, N346, N378, N95);
  xnor KeyGate_0_112(KeyNOTWire_0[48], keyIn_0_112, KeyWire_0[112]);
  not KeyNOTGate_0_48(N411, KeyNOTWire_0[48]);
  nand NAND4_146 (KeyWire_0[113], N259, N347, N379, N108);
  xnor KeyGate_0_113(KeyNOTWire_0[49], keyIn_0_113, KeyWire_0[113]);
  not KeyNOTGate_0_49(N414, KeyNOTWire_0[49]);
  not NOT1_147 (KeyWire_0[114], N380);
  xnor KeyGate_0_114(KeyNOTWire_0[50], keyIn_0_114, KeyWire_0[114]);
  not KeyNOTGate_0_50(N415, KeyNOTWire_0[50]);
  and AND8_148 (KeyWire_0[115], N381, N386, N393, N399, N404, N407, N411, N414);
  xor KeyGate_0_115(N416, keyIn_0_115, KeyWire_0[115]);
  not NOT1_149 (KeyWire_0[116], N393);
  xor KeyGate_0_116(N417, keyIn_0_116, KeyWire_0[116]);
  not NOT1_150 (KeyWire_0[117], N404);
  xor KeyGate_0_117(N418, keyIn_0_117, KeyWire_0[117]);
  not NOT1_151 (KeyWire_0[118], N407);
  xnor KeyGate_0_118(N419, keyIn_0_118, KeyWire_0[118]);
  not NOT1_152 (KeyWire_0[119], N411);
  xnor KeyGate_0_119(KeyNOTWire_0[51], keyIn_0_119, KeyWire_0[119]);
  not KeyNOTGate_0_51(N420, KeyNOTWire_0[51]);
  nor NOR2_153 (KeyWire_0[120], N415, N416);
  xnor KeyGate_0_120(KeyNOTWire_0[52], keyIn_0_120, KeyWire_0[120]);
  not KeyNOTGate_0_52(N421, KeyNOTWire_0[52]);
  nand NAND2_154 (KeyWire_0[121], N386, N417);
  xnor KeyGate_0_121(N422, keyIn_0_121, KeyWire_0[121]);
  nand NAND4_155 (KeyWire_0[122], N386, N393, N418, N399);
  xor KeyGate_0_122(KeyNOTWire_0[53], keyIn_0_122, KeyWire_0[122]);
  not KeyNOTGate_0_53(N425, KeyNOTWire_0[53]);
  nand NAND3_156 (KeyWire_0[123], N399, N393, N419);
  xor KeyGate_0_123(N428, keyIn_0_123, KeyWire_0[123]);
  nand NAND4_157 (KeyWire_0[124], N386, N393, N407, N420);
  xnor KeyGate_0_124(KeyNOTWire_0[54], keyIn_0_124, KeyWire_0[124]);
  not KeyNOTGate_0_54(N429, KeyNOTWire_0[54]);
  nand NAND4_158 (KeyWire_0[125], N381, N386, N422, N399);
  xnor KeyGate_0_125(KeyNOTWire_0[55], keyIn_0_125, KeyWire_0[125]);
  not KeyNOTGate_0_55(N430, KeyNOTWire_0[55]);
  nand NAND4_159 (KeyWire_0[126], N381, N386, N425, N428);
  xor KeyGate_0_126(KeyNOTWire_0[56], keyIn_0_126, KeyWire_0[126]);
  not KeyNOTGate_0_56(N431, KeyNOTWire_0[56]);
  nand NAND4_160 (KeyWire_0[127], N381, N422, N425, N429);
  xnor KeyGate_0_127(N432, keyIn_0_127, KeyWire_0[127]);

endmodule
