// Verilog File 
module top (G101,G104,G107,G110,G113,G116,G119,G122,G125,
G128,G131,G134,G137,G140,G143,G146,G210,G214,G217,
G221,G224,G227,G234,G237,G469,G472,G475,G478,G898,
G900,G902,G952,G953,G3,G6,G9,G12,G30,G45,
G48,G15,G18,G21,G24,G27,G33,G36,G39,G42,
G75,G51,G54,G60,G63,G66,G69,G72,G57,keyinput0,
keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,
keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,
keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,
keyinput31,keyinput32,keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,
keyinput41,keyinput42,keyinput43,keyinput44,keyinput45,keyinput46,keyinput47);

input G101,G104,G107,G110,G113,G116,G119,G122,G125,
G128,G131,G134,G137,G140,G143,G146,G210,G214,G217,
G221,G224,G227,G234,G237,G469,G472,G475,G478,G898,
G900,G902,G952,G953,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,
keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,
keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,
keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,keyinput35,
keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,keyinput45,
keyinput46,keyinput47;

output G3,G6,G9,G12,G30,G45,G48,G15,G18,
G21,G24,G27,G33,G36,G39,G42,G75,G51,G54,
G60,G63,G66,G69,G72,G57;

wire G149,G153,G156,G160,G165,G168,G171,G175,G179,
G184,G188,G191,G194,G198,G202,G206,G231,G233,G241,
G244,G245,G248,G517,G529,G541,G553,G859,G862,G907,
G909,G911,G918,G919,G922,G926,G930,G932,G934,G938,
G943,G947,G949,G1506,G1514,G1522,G1530,G1538,G1546,G1554,
G1562,G1570,G1578,G1586,G1594,G1602,G1610,G1618,G1626,G1512,
G1520,G1528,G1536,G1544,G1552,G1560,G1568,G1576,G1584,G1592,
G1600,G1608,G1616,G1624,G1632,G50,G52,G56,G58,G62,
G64,G251,G254,G288,G291,G299,G302,G318,G321,G327,
G330,G352,G355,G369,G382,G385,G853,G856,G893,G954,
G955,G1050,G1053,G1176,G1179,G1197,G1207,G1222,G1244,G1278,
G1290,G1300,G1312,G1332,G1335,G1442,G1450,G1458,G1466,G1474,
G1482,G1490,G1498,G1634,G1644,G1657,G1665,G1697,G1705,G1713,
G1721,G1745,G1753,G1785,G1793,G1814,G1817,G1830,G1833,G1841,
G1849,G1854,G1857,G1870,G1873,G1878,G1881,G1642,G1652,G1056,
G1057,G1182,G1183,G1211,G1298,G1320,G1338,G1339,G457,G459,
G482,G487,G492,G505,G1456,G1448,G1472,G1464,G1488,G1480,
G1504,G1496,G956,G967,G978,G979,G980,G1661,G990,G1669,
G1030,G1701,G1040,G1709,G1058,G1717,G1068,G1725,G1078,G1090,
G1100,G1749,G1112,G1757,G1154,G1789,G1166,G1797,G1194,G1201,
G1204,G1820,G1821,G1230,G1836,G1837,G1252,G1256,G1845,G1268,
G1853,G1860,G1861,G1286,G1876,G1877,G1308,G1884,G1885,G1654,
G1662,G1694,G1702,G1710,G1718,G1726,G1734,G1742,G1750,G1782,
G1790,G1838,G1846,G297,G298,G361,G362,G404,G405,G1225,
G1226,G1247,G1248,G1281,G1282,G1303,G1304,G1315,G1316,G998,
G988,G268,G1038,G1048,G1076,G1066,G1098,G1120,G1174,G363,
G1210,G373,G1276,G406,G565,G566,G614,G615,G958,G969,
G1660,G984,G1668,G994,G1700,G1034,G1708,G1044,G1716,G1062,
G1724,G1072,G1732,G1086,G1740,G1748,G1104,G1108,G1756,G1116,
G1788,G1158,G1162,G1796,G1170,G1200,G1203,G1227,G1249,G1844,
G1260,G1264,G1852,G1272,G1283,G1305,G1317,G1410,G1418,G1426,
G1434,G269,G372,G983,G993,G1033,G1043,G1061,G1071,G1103,
G1115,G1157,G1169,G1184,G1202,G1259,G1271,G1322,G374,G396,
G1321,G1424,G1416,G1440,G1432,G985,G995,G1035,G1045,G1063,
G1073,G1105,G1117,G1159,G1171,G1212,G1231,G1232,G1253,G1254,
G1261,G1273,G1287,G1288,G1309,G1310,G1192,G397,G1330,G1000,
G1010,G1233,G1255,G1289,G1311,G1381,G257,G999,G260,G989,
G272,G1039,G294,G1049,G305,G1077,G308,G1067,G333,G1121,
G358,G1175,G1220,G388,G1277,G398,G1109,G1110,G1163,G1164,
G1234,G1265,G1266,G1822,G1862,G1865,G258,G261,G273,G1018,
G1008,G295,G306,G309,G334,G359,G389,G1385,G1111,G1165,
G1267,G1886,G259,G262,G274,G296,G307,G310,G335,G360,
G1242,G390,G1828,G1868,G1869,G1373,G1798,G1825,G265,G314,
G336,G407,G1293,G1294,G1892,G1777,G1889,G410,G1377,G1804,
G1237,G1829,G1295,G1670,G1678,G1729,G1737,G1761,G1769,G340,
G343,G1781,G1238,G1325,G1893,G1340,G1352,G1673,G1681,G1801,
G1897,G1905,G391,G1299,G1676,G1684,G1081,G1733,G1093,G1741,
G1765,G1773,G1239,G1326,G1894,G1902,G392,G1360,G1003,G1677,
G1013,G1685,G1082,G1094,G1122,G1134,G1187,G1805,G1327,G1901,
G1348,G1909,G1758,G1766,G377,G1243,G393,G1004,G1014,G1083,
G1095,G1188,G1900,G1344,G1908,G1356,G1142,G378,G399,G1331,
G1005,G1015,G1764,G1126,G1130,G1772,G1138,G1189,G1343,G1355,
G324,G1099,G379,G400,G449,G1087,G1088,G1125,G1137,G1345,
G1357,G1397,G277,G1019,G280,G1009,G325,G364,G1193,G401,
G1089,G1127,G1139,G278,G281,G326,G365,G413,G1361,G1401,
G445,G1349,G1350,G1389,G1493,G1501,G1689,G279,G282,G346,
G1143,G366,G414,G453,G1131,G1132,G1351,G1365,G1405,G285,
G347,G367,G415,G1393,G556,G1505,G559,G1497,G1693,G1133,
G1477,G1485,G1809,G348,G1369,G1409,G557,G560,G1362,G1378,
G1429,G1437,G1686,G1774,G1910,G1918,G544,G1489,G547,G1481,
G558,G561,G1813,G1370,G1368,G417,G1384,G424,G508,G1441,
G511,G1433,G545,G548,G564,G1692,G1024,G1780,G1148,G1916,
G1924,G416,G1376,G421,G423,G509,G512,G546,G549,G719,
G722,G1023,G1147,G418,G420,G425,G510,G513,G552,G1025,
G1149,G419,G422,G441,G516,G725,G728,G1029,G1153,G433,
G437,G663,G666,G731,G746,G756,G770,G1461,G1469,G1413,
G1421,G1445,G1453,G532,G1473,G535,G1465,G495,G1425,G498,
G1417,G520,G1457,G523,G1449,G533,G536,G496,G499,G521,
G524,G534,G537,G497,G500,G522,G525,G540,G503,G528,
G669,G672,G569,G588,G618,G639,G867,G588a,G588b,G639a,
G639b,G675,G688,G696,G710,G73,G572,G573,G621,G622,
G776,G780,G784,G788,G812,G832,G836,G1509,G1517,G1525,
G1533,G1581,G1621,G1629,G792,G796,G800,G804,G808,G816,
G820,G824,G828,G871,G873,G875,G877,G879,G881,G883,
G885,G1541,G1549,G1557,G1565,G1573,G1589,G1597,G1605,G1613,
G1,G1513,G4,G1521,G7,G1529,G10,G1537,G28,G1585,
G43,G1625,G46,G1633,G886,G2,G5,G8,G11,G13,
G1545,G16,G1553,G19,G1561,G22,G1569,G25,G1577,G29,
G31,G1593,G34,G1601,G37,G1609,G40,G1617,G44,G47,
G857,G860,G863,G865,G14,G17,G20,G23,G26,G32,
G35,G38,G41,G1913,G1921,G887,G462,G74,G1637,G1917,
G1647,G1925,G1020,G1144,G1386,G1394,G1402,G1638,G1648,G1806,
G1639,G1649,G287,G350,G427,G429,G431,G1028,G1152,G1392,
G1400,G1408,G1812,G1216,G286,G349,G426,G428,G430,G67,
G1643,G70,G1653,G1215,G49,G53,G59,G61,G65,G68,
G71,G1217,G375,G1221,G376,G55,muxed0,muxed1,muxed2,muxed3,
muxed4,muxed5,muxed6,muxed7,muxed8,muxed9,muxed10,muxed11,muxed12,muxed13,
muxed14,muxed15,muxed16,muxed17,muxed18,muxed19,muxed20,muxed21,muxed22,muxed23,
muxed24,muxed25,muxed26,muxed27,muxed28,muxed29,muxed30,muxed31,muxed32,muxed33,
muxed34,muxed35,muxed36,muxed37,muxed38,muxed39,muxed40,muxed41,muxed42,muxed43,
muxed44,muxed45,muxed46,muxed47;
not gate_0(G149,G101);
not gate_1(G153,G104);
not gate_2(G156,G107);
not gate_3(G160,G110);
not gate_4(G165,G113);
not gate_5(G168,G116);
not gate_6(G171,G119);
not gate_7(G175,G122);
not gate_8(G179,G125);
not gate_9(G184,G128);
not gate_10(G188,G131);
not gate_11(G191,G134);
not gate_12(G194,G137);
not gate_13(G198,G140);
not gate_14(G202,G143);
not gate_15(G206,G146);
nand gate_16(G231,G224,G898);
nand gate_17(G233,G227,G900);
not gate_18(G241,G237);
not gate_19(G244,G237);
buf gate_20(G245,G234);
buf gate_21(G248,G234);
not gate_22(G517,G469);
not gate_23(G529,G472);
not gate_24(G541,G475);
not gate_25(G553,G478);
not gate_26(G859,G953);
not gate_27(G862,G953);
not gate_28(G907,G898);
not gate_29(G909,G900);
buf gate_30(G911,G902);
not gate_31(G918,G902);
buf gate_32(G919,G902);
not gate_33(G922,G902);
buf gate_34(G926,G952);
not gate_35(G930,G952);
not gate_36(G932,G952);
buf gate_37(G934,G953);
not gate_38(G938,G953);
buf gate_39(G943,G953);
buf gate_40(G947,G953);
not gate_41(G949,G953);
buf gate_42(G1506,G101);
buf gate_43(G1514,G104);
buf gate_44(G1522,G107);
buf gate_45(G1530,G110);
buf gate_46(G1538,G113);
buf gate_47(G1546,G116);
buf gate_48(G1554,G119);
buf gate_49(G1562,G122);
buf gate_50(G1570,G125);
buf gate_51(G1578,G128);
buf gate_52(G1586,G131);
buf gate_53(G1594,G134);
buf gate_54(G1602,G137);
buf gate_55(G1610,G140);
buf gate_56(G1618,G143);
buf gate_57(G1626,G146);
not gate_58(G1512,G1506);
not gate_59(G1520,G1514);
not gate_60(G1528,G1522);
not gate_61(G1536,G1530);
not gate_62(G1544,G1538);
not gate_63(G1552,G1546);
not gate_64(G1560,G1554);
not gate_65(G1568,G1562);
not gate_66(G1576,G1570);
not gate_67(G1584,G1578);
not gate_68(G1592,G1586);
not gate_69(G1600,G1594);
not gate_70(G1608,G1602);
not gate_71(G1616,G1610);
not gate_72(G1624,G1618);
not gate_73(G1632,G1626);
nand gate_74(G50,G930,G947);
nand gate_75(G52,G930,G947);
nand gate_76(G56,G930,G947);
nand gate_77(G58,G930,G947);
nand gate_78(G62,G930,G947);
nand gate_79(G64,G930,G947);
buf gate_80(G251,G149);
buf gate_81(G254,G153);
buf gate_82(G288,G165);
buf gate_83(G291,G168);
buf gate_84(G299,G184);
buf gate_85(G302,G202);
and gate_86(G318,G224,G938);
buf gate_87(G321,G179);
buf gate_88(G327,G188);
buf gate_89(G330,G191);
and gate_90(G352,G227,G938);
buf gate_91(G355,G198);
and gate_92(G369,G210,G241,G938);
buf gate_93(G382,G206);
buf gate_94(G385,G198);
nand gate_95(G853,G943,G907);
nand gate_96(G856,G943,G909);
nand gate_97(G893,G248,G237);
nand gate_98(G954,G248,G922);
nand gate_99(G955,G244,G922);
buf gate_100(G1050,G160);
buf gate_101(G1053,G175);
buf gate_102(G1176,G179);
buf gate_103(G1179,G198);
buf gate_104(G1197,G149);
buf gate_105(G1207,G149);
buf gate_106(G1222,G153);
buf gate_107(G1244,G188);
buf gate_108(G1278,G156);
and gate_109(G1290,G217,G245,G938);
buf gate_110(G1300,G191);
buf gate_111(G1312,G160);
buf gate_112(G1332,G194);
and gate_113(G1335,G221,G245,G938);
buf gate_114(G1442,G517);
buf gate_115(G1450,G517);
buf gate_116(G1458,G529);
buf gate_117(G1466,G529);
buf gate_118(G1474,G541);
buf gate_119(G1482,G541);
buf gate_120(G1490,G553);
buf gate_121(G1498,G553);
and gate_122(G1634,G231,G934);
and gate_123(G1644,G233,G934);
buf gate_124(G1657,G156);
buf gate_125(G1665,G156);
buf gate_126(G1697,G171);
buf gate_127(G1705,G171);
buf gate_128(G1713,G206);
buf gate_129(G1721,G206);
buf gate_130(G1745,G194);
buf gate_131(G1753,G194);
buf gate_132(G1785,G160);
buf gate_133(G1793,G160);
buf gate_134(G1814,G165);
buf gate_135(G1817,G175);
and gate_136(G1830,G214,G241,G938);
buf gate_137(G1833,G202);
buf gate_138(G1841,G179);
buf gate_139(G1849,G179);
buf gate_140(G1854,G168);
buf gate_141(G1857,G175);
buf gate_142(G1870,G184);
buf gate_143(G1873,G202);
buf gate_144(G1878,G171);
buf gate_145(G1881,G184);
not gate_146(G1642,G1634);
not gate_147(G1652,G1644);
not gate_148(G1056,muxed24);
not gate_149(G1057,G1053);
not gate_150(G1182,G1176);
not gate_151(G1183,G1179);
not gate_152(G1211,G1207);
not gate_153(G1298,G1290);
not gate_154(G1320,G1312);
not gate_155(G1338,G1332);
not gate_156(G1339,G1335);
and gate_157(G457,G210,G955);
and gate_158(G459,G217,G954);
nand gate_159(G482,G214,G955);
nand gate_160(G487,G221,G954);
nand gate_161(G492,G210,G955);
nand gate_162(G505,G217,G954);
not gate_163(G1456,G1450);
not gate_164(G1448,G1442);
not gate_165(G1472,G1466);
not gate_166(G1464,G1458);
not gate_167(G1488,G1482);
not gate_168(G1480,G1474);
not gate_169(G1504,G1498);
not gate_170(G1496,G1490);
nand gate_171(G956,G907,G919,G943,G893);
nand gate_172(G967,G909,G919,G943,G893);
nand gate_173(G978,G926,G949,G893);
and gate_174(G979,G926,G949,G893);
buf gate_175(G980,G251);
not gate_176(G1661,G1657);
buf gate_177(G990,G251);
not gate_178(G1669,G1665);
buf gate_179(G1030,G288);
not gate_180(G1701,G1697);
buf gate_181(G1040,G288);
not gate_182(G1709,G1705);
buf gate_183(G1058,G299);
not gate_184(G1717,G1713);
buf gate_185(G1068,G299);
not gate_186(G1725,G1721);
buf gate_187(G1078,G318);
buf gate_188(G1090,G318);
buf gate_189(G1100,G327);
not gate_190(G1749,G1745);
buf gate_191(G1112,G327);
not gate_192(G1757,G1753);
buf gate_193(G1154,G352);
not gate_194(G1789,G1785);
buf gate_195(G1166,G352);
not gate_196(G1797,G1793);
buf gate_197(G1194,G369);
not gate_198(G1201,G1197);
buf gate_199(G1204,G369);
not gate_200(G1820,G1814);
not gate_201(G1821,G1817);
not gate_202(G1230,G1222);
not gate_203(G1836,G1830);
not gate_204(G1837,G1833);
not gate_205(G1252,G1244);
buf gate_206(G1256,G382);
not gate_207(G1845,G1841);
buf gate_208(G1268,G382);
not gate_209(G1853,G1849);
not gate_210(G1860,G1854);
not gate_211(G1861,G1857);
not gate_212(G1286,G1278);
not gate_213(G1876,G1870);
not gate_214(G1877,G1873);
not gate_215(G1308,G1300);
not gate_216(G1884,G1878);
not gate_217(G1885,G1881);
buf gate_218(G1654,G254);
buf gate_219(G1662,G254);
buf gate_220(G1694,G291);
buf gate_221(G1702,G291);
buf gate_222(G1710,G302);
buf gate_223(G1718,G302);
buf gate_224(G1726,G321);
buf gate_225(G1734,G321);
buf gate_226(G1742,G330);
buf gate_227(G1750,G330);
buf gate_228(G1782,G355);
buf gate_229(G1790,G355);
buf gate_230(G1838,G385);
buf gate_231(G1846,G385);
nand gate_232(G297,G1053,G1056);
nand gate_233(G298,muxed24,G1057);
nand gate_234(G361,G1179,G1182);
nand gate_235(G362,G1176,G1183);
nand gate_236(G404,G1335,G1338);
nand gate_237(G405,G1332,G1339);
nand gate_238(G1225,G1817,G1820);
nand gate_239(G1226,G1814,G1821);
nand gate_240(G1247,G1833,G1836);
nand gate_241(G1248,G1830,G1837);
nand gate_242(G1281,G1857,G1860);
nand gate_243(G1282,G1854,G1861);
nand gate_244(G1303,G1873,G1876);
nand gate_245(G1304,G1870,G1877);
nand gate_246(G1315,G1881,G1884);
nand gate_247(G1316,G1878,G1885);
not gate_248(G998,muxed12);
not gate_249(G988,G980);
nand gate_250(G268,G297,G298);
not gate_251(G1038,G1030);
not gate_252(G1048,G1040);
not gate_253(G1076,G1068);
not gate_254(G1066,G1058);
not gate_255(G1098,G1090);
not gate_256(G1120,G1112);
not gate_257(G1174,G1166);
nand gate_258(G363,G361,G362);
not gate_259(G1210,G1204);
nand gate_260(G373,G1204,G1211);
not gate_261(G1276,G1268);
nand gate_262(G406,G404,G405);
not gate_263(G565,G482);
buf gate_264(G566,G482);
not gate_265(G614,G487);
buf gate_266(G615,G487);
nand gate_267(G958,G956,G978);
nand gate_268(G969,G967,G978);
not gate_269(G1660,G1654);
nand gate_270(G984,G1654,G1661);
not gate_271(G1668,G1662);
nand gate_272(G994,G1662,G1669);
not gate_273(G1700,G1694);
nand gate_274(G1034,G1694,G1701);
not gate_275(G1708,G1702);
nand gate_276(G1044,G1702,G1709);
not gate_277(G1716,G1710);
nand gate_278(G1062,G1710,G1717);
not gate_279(G1724,G1718);
nand gate_280(G1072,G1718,G1725);
not gate_281(G1732,G1726);
not gate_282(G1086,G1078);
not gate_283(G1740,G1734);
not gate_284(G1748,G1742);
nand gate_285(G1104,G1742,G1749);
not gate_286(G1108,G1100);
not gate_287(G1756,G1750);
nand gate_288(G1116,G1750,G1757);
not gate_289(G1788,G1782);
nand gate_290(G1158,G1782,G1789);
not gate_291(G1162,G1154);
not gate_292(G1796,G1790);
nand gate_293(G1170,G1790,G1797);
not gate_294(G1200,G1194);
nand gate_295(G1203,G1194,G1201);
nand gate_296(G1227,G1225,G1226);
nand gate_297(G1249,G1247,G1248);
not gate_298(G1844,G1838);
nand gate_299(G1260,G1838,G1845);
not gate_300(G1264,G1256);
not gate_301(G1852,G1846);
nand gate_302(G1272,G1846,G1853);
nand gate_303(G1283,G1281,G1282);
nand gate_304(G1305,G1303,G1304);
nand gate_305(G1317,G1315,G1316);
buf gate_306(G1410,G492);
buf gate_307(G1418,G492);
buf gate_308(G1426,G505);
buf gate_309(G1434,G505);
not gate_310(G269,G268);
nand gate_311(G372,G1207,G1210);
nand gate_312(G983,G1657,G1660);
nand gate_313(G993,G1665,G1668);
nand gate_314(G1033,G1697,G1700);
nand gate_315(G1043,G1705,G1708);
nand gate_316(G1061,G1713,G1716);
nand gate_317(G1071,G1721,G1724);
nand gate_318(G1103,G1745,G1748);
nand gate_319(G1115,G1753,G1756);
nand gate_320(G1157,G1785,G1788);
nand gate_321(G1169,G1793,G1796);
not gate_322(G1184,G363);
nand gate_323(G1202,G1197,G1200);
nand gate_324(G1259,G1841,G1844);
nand gate_325(G1271,G1849,G1852);
not gate_326(G1322,G406);
nand gate_327(G374,G372,G373);
nand gate_328(G396,G1317,G1320);
not gate_329(G1321,G1317);
not gate_330(G1424,G1418);
not gate_331(G1416,G1410);
not gate_332(G1440,G1434);
not gate_333(G1432,G1426);
nand gate_334(G985,muxed0,G984);
nand gate_335(G995,G993,G994);
nand gate_336(G1035,G1033,G1034);
nand gate_337(G1045,G1043,G1044);
nand gate_338(G1063,G1061,G1062);
nand gate_339(G1073,G1071,G1072);
nand gate_340(G1105,G1103,G1104);
nand gate_341(G1117,G1115,G1116);
nand gate_342(G1159,G1157,G1158);
nand gate_343(G1171,G1169,G1170);
nand gate_344(G1212,G1202,G1203);
not gate_345(G1231,G1227);
nand gate_346(G1232,G1227,G1230);
not gate_347(G1253,G1249);
nand gate_348(G1254,G1249,G1252);
nand gate_349(G1261,G1259,G1260);
nand gate_350(G1273,G1271,G1272);
not gate_351(G1287,G1283);
nand gate_352(G1288,G1283,G1286);
not gate_353(G1309,G1305);
nand gate_354(G1310,G1305,G1308);
not gate_355(G1192,muxed8);
nand gate_356(G397,G1312,G1321);
not gate_357(G1330,G1322);
buf gate_358(G1000,G269);
buf gate_359(G1010,G269);
nand gate_360(G1233,G1222,G1231);
nand gate_361(G1255,G1244,G1253);
nand gate_362(G1289,G1278,G1287);
nand gate_363(G1311,G1300,G1309);
not gate_364(G1381,G374);
nand gate_365(G257,G995,G998);
not gate_366(G999,G995);
nand gate_367(G260,muxed11,G988);
not gate_368(G989,muxed11);
nand gate_369(G272,G1035,G1038);
not gate_370(G1039,G1035);
nand gate_371(G294,G1045,G1048);
not gate_372(G1049,G1045);
nand gate_373(G305,G1073,G1076);
not gate_374(G1077,G1073);
nand gate_375(G308,G1063,G1066);
not gate_376(G1067,G1063);
nand gate_377(G333,G1117,G1120);
not gate_378(G1121,G1117);
nand gate_379(G358,G1171,G1174);
not gate_380(G1175,G1171);
not gate_381(G1220,G1212);
nand gate_382(G388,G1273,G1276);
not gate_383(G1277,G1273);
nand gate_384(G398,G396,G397);
not gate_385(G1109,G1105);
nand gate_386(G1110,G1105,G1108);
not gate_387(G1163,G1159);
nand gate_388(G1164,G1159,G1162);
nand gate_389(G1234,G1232,G1233);
not gate_390(G1265,G1261);
nand gate_391(G1266,G1261,G1264);
nand gate_392(G1822,G1254,G1255);
nand gate_393(G1862,G1310,G1311);
nand gate_394(G1865,G1288,G1289);
nand gate_395(G258,muxed12,G999);
nand gate_396(G261,G980,muxed9);
nand gate_397(G273,G1030,G1039);
not gate_398(G1018,G1010);
not gate_399(G1008,G1000);
nand gate_400(G295,G1040,G1049);
nand gate_401(G306,G1068,G1077);
nand gate_402(G309,G1058,G1067);
nand gate_403(G334,G1112,G1121);
nand gate_404(G359,G1166,G1175);
nand gate_405(G389,G1268,G1277);
not gate_406(G1385,G1381);
nand gate_407(G1111,G1100,G1109);
nand gate_408(G1165,G1154,G1163);
nand gate_409(G1267,G1256,muxed44);
not gate_410(G1886,G398);
nand gate_411(G259,G257,muxed23);
nand gate_412(G262,G260,muxed7);
nand gate_413(G274,G272,G273);
nand gate_414(G296,G294,G295);
nand gate_415(G307,G305,G306);
nand gate_416(G310,G308,G309);
nand gate_417(G335,G333,G334);
nand gate_418(G360,G358,G359);
not gate_419(G1242,G1234);
nand gate_420(G390,G388,G389);
not gate_421(G1828,G1822);
not gate_422(G1868,G1862);
not gate_423(G1869,G1865);
nand gate_424(G1373,G1164,G1165);
nand gate_425(G1798,G1110,G1111);
nand gate_426(G1825,G1266,G1267);
not gate_427(G265,muxed21);
not gate_428(G314,G307);
not gate_429(G336,G335);
not gate_430(G407,G296);
nand gate_431(G1293,G1865,G1868);
nand gate_432(G1294,G1862,G1869);
not gate_433(G1892,muxed18);
not gate_434(G1777,G360);
not gate_435(G1889,G390);
buf gate_436(G410,G310);
not gate_437(G1377,G1373);
not gate_438(G1804,G1798);
nand gate_439(G1237,G1825,G1828);
not gate_440(G1829,G1825);
nand gate_441(G1295,G1293,G1294);
buf gate_442(G1670,G274);
buf gate_443(G1678,G274);
buf gate_444(G1729,G310);
buf gate_445(G1737,G310);
buf gate_446(G1761,muxed6);
buf gate_447(G1769,muxed6);
buf gate_448(G340,G336);
buf gate_449(G343,muxed36);
not gate_450(G1781,G1777);
nand gate_451(G1238,G1822,G1829);
nand gate_452(G1325,G1889,G1892);
not gate_453(G1893,G1889);
buf gate_454(G1340,G407);
buf gate_455(G1352,G407);
buf gate_456(G1673,muxed20);
buf gate_457(G1681,muxed20);
buf gate_458(G1801,muxed36);
buf gate_459(G1897,G336);
buf gate_460(G1905,G336);
nand gate_461(G391,G1295,G1298);
not gate_462(G1299,G1295);
not gate_463(G1676,G1670);
not gate_464(G1684,G1678);
nand gate_465(G1081,G1729,G1732);
not gate_466(G1733,G1729);
nand gate_467(G1093,G1737,G1740);
not gate_468(G1741,G1737);
not gate_469(G1765,G1761);
not gate_470(G1773,muxed5);
nand gate_471(G1239,G1237,G1238);
nand gate_472(G1326,muxed18,G1893);
buf gate_473(G1894,G410);
buf gate_474(G1902,G410);
nand gate_475(G392,G1290,G1299);
not gate_476(G1360,G1352);
nand gate_477(G1003,G1673,G1676);
not gate_478(G1677,G1673);
nand gate_479(G1013,muxed19,G1684);
not gate_480(G1685,muxed19);
nand gate_481(G1082,G1726,G1733);
nand gate_482(G1094,G1734,G1741);
buf gate_483(G1122,G340);
buf gate_484(G1134,G340);
nand gate_485(G1187,G1801,G1804);
not gate_486(G1805,G1801);
nand gate_487(G1327,G1325,G1326);
not gate_488(G1901,G1897);
not gate_489(G1348,G1340);
not gate_490(G1909,G1905);
buf gate_491(G1758,G343);
buf gate_492(G1766,G343);
nand gate_493(G377,G1239,G1242);
not gate_494(G1243,G1239);
nand gate_495(G393,G391,G392);
nand gate_496(G1004,G1670,G1677);
nand gate_497(G1014,G1678,muxed17);
nand gate_498(G1083,G1081,G1082);
nand gate_499(G1095,G1093,G1094);
nand gate_500(G1188,G1798,G1805);
not gate_501(G1900,G1894);
nand gate_502(G1344,G1894,G1901);
not gate_503(G1908,G1902);
nand gate_504(G1356,G1902,G1909);
not gate_505(G1142,G1134);
nand gate_506(G378,G1234,G1243);
nand gate_507(G399,G1327,G1330);
not gate_508(G1331,G1327);
nand gate_509(G1005,G1003,G1004);
nand gate_510(G1015,G1013,muxed15);
not gate_511(G1764,G1758);
nand gate_512(G1126,G1758,G1765);
not gate_513(G1130,G1122);
not gate_514(G1772,G1766);
nand gate_515(G1138,G1766,G1773);
nand gate_516(G1189,G1187,G1188);
nand gate_517(G1343,G1897,G1900);
nand gate_518(G1355,G1905,G1908);
nand gate_519(G324,G1095,G1098);
not gate_520(G1099,G1095);
nand gate_521(G379,G377,G378);
nand gate_522(G400,G1322,G1331);
nand gate_523(G449,G393,G918);
not gate_524(G1087,G1083);
nand gate_525(G1088,G1083,G1086);
nand gate_526(G1125,G1761,G1764);
nand gate_527(G1137,muxed5,G1772);
nand gate_528(G1345,G1343,G1344);
nand gate_529(G1357,G1355,G1356);
buf gate_530(G1397,G393);
nand gate_531(G277,muxed14,G1018);
not gate_532(G1019,muxed14);
nand gate_533(G280,G1005,G1008);
not gate_534(G1009,G1005);
nand gate_535(G325,G1090,G1099);
nand gate_536(G364,G1189,G1192);
not gate_537(G1193,G1189);
nand gate_538(G401,G399,G400);
nand gate_539(G1089,G1078,G1087);
nand gate_540(G1127,G1125,G1126);
nand gate_541(G1139,muxed3,G1138);
nand gate_542(G278,G1010,muxed13);
nand gate_543(G281,G1000,G1009);
nand gate_544(G326,G324,G325);
nand gate_545(G365,muxed8,G1193);
nand gate_546(G413,G1357,G1360);
not gate_547(G1361,G1357);
not gate_548(G1401,G1397);
nand gate_549(G445,G379,G918);
not gate_550(G1349,G1345);
nand gate_551(G1350,G1345,G1348);
buf gate_552(G1389,G379);
buf gate_553(G1493,muxed37);
buf gate_554(G1501,muxed37);
nand gate_555(G1689,G1088,G1089);
nand gate_556(G279,G277,G278);
nand gate_557(G282,G280,G281);
nand gate_558(G346,muxed2,G1142);
not gate_559(G1143,muxed2);
nand gate_560(G366,G364,G365);
nand gate_561(G414,G1352,G1361);
nand gate_562(G453,G401,G918);
not gate_563(G1131,G1127);
nand gate_564(G1132,G1127,G1130);
nand gate_565(G1351,G1340,G1349);
not gate_566(G1365,G326);
buf gate_567(G1405,G401);
not gate_568(G285,G279);
nand gate_569(G347,G1134,muxed1);
not gate_570(G367,G366);
nand gate_571(G415,G413,G414);
not gate_572(G1393,G1389);
nand gate_573(G556,G1501,G1504);
not gate_574(G1505,G1501);
nand gate_575(G559,muxed47,G1496);
not gate_576(G1497,muxed47);
not gate_577(G1693,G1689);
nand gate_578(G1133,G1122,G1131);
buf gate_579(G1477,G445);
buf gate_580(G1485,G445);
nand gate_581(G1809,G1350,G1351);
nand gate_582(G348,G346,G347);
not gate_583(G1369,G1365);
not gate_584(G1409,G1405);
nand gate_585(G557,G1498,G1505);
nand gate_586(G560,G1490,muxed45);
buf gate_587(G1362,G282);
not gate_588(G1378,G415);
buf gate_589(G1429,G453);
buf gate_590(G1437,G453);
buf gate_591(G1686,G282);
nand gate_592(G1774,G1132,G1133);
and gate_593(G1910,G285,G853);
and gate_594(G1918,G856,G367);
nand gate_595(G544,G1485,G1488);
not gate_596(G1489,G1485);
nand gate_597(G547,G1477,G1480);
not gate_598(G1481,G1477);
nand gate_599(G558,G556,G557);
nand gate_600(G561,G559,muxed43);
not gate_601(G1813,G1809);
not gate_602(G1370,G348);
not gate_603(G1368,G1362);
nand gate_604(G417,G1362,G1369);
not gate_605(G1384,G1378);
nand gate_606(G424,G1378,G1385);
nand gate_607(G508,G1437,G1440);
not gate_608(G1441,G1437);
nand gate_609(G511,G1429,G1432);
not gate_610(G1433,G1429);
nand gate_611(G545,G1482,G1489);
nand gate_612(G548,G1474,G1481);
not gate_613(G564,G558);
not gate_614(G1692,G1686);
nand gate_615(G1024,G1686,G1693);
not gate_616(G1780,G1774);
nand gate_617(G1148,G1774,G1781);
not gate_618(G1916,G1910);
not gate_619(G1924,G1918);
nand gate_620(G416,G1365,G1368);
not gate_621(G1376,G1370);
nand gate_622(G421,G1370,G1377);
nand gate_623(G423,G1381,G1384);
nand gate_624(G509,G1434,G1441);
nand gate_625(G512,G1426,G1433);
nand gate_626(G546,G544,G545);
nand gate_627(G549,G547,G548);
not gate_628(G719,muxed42);
buf gate_629(G722,muxed42);
nand gate_630(G1023,G1689,G1692);
nand gate_631(G1147,G1777,G1780);
nand gate_632(G418,G416,G417);
nand gate_633(G420,G1373,G1376);
nand gate_634(G425,G423,G424);
nand gate_635(G510,G508,G509);
nand gate_636(G513,G511,G512);
not gate_637(G552,G546);
nand gate_638(G1025,G1023,G1024);
nand gate_639(G1149,G1147,G1148);
not gate_640(G419,G418);
nand gate_641(G422,G420,G421);
nand gate_642(G441,G425,G918);
not gate_643(G516,G510);
not gate_644(G725,muxed34);
buf gate_645(G728,muxed34);
not gate_646(G1029,G1025);
not gate_647(G1153,G1149);
nand gate_648(G433,G419,G918);
nand gate_649(G437,G422,G918);
not gate_650(G663,G513);
buf gate_651(G666,G513);
and gate_652(G731,G719,G725);
and gate_653(G746,muxed41,G725);
and gate_654(G756,G719,G728);
and gate_655(G770,muxed41,G728);
buf gate_656(G1461,G441);
buf gate_657(G1469,G441);
buf gate_658(G1413,G433);
buf gate_659(G1421,G433);
buf gate_660(G1445,G437);
buf gate_661(G1453,G437);
nand gate_662(G532,G1469,G1472);
not gate_663(G1473,G1469);
nand gate_664(G535,muxed25,G1464);
not gate_665(G1465,muxed25);
nand gate_666(G495,G1421,G1424);
not gate_667(G1425,G1421);
nand gate_668(G498,G1413,G1416);
not gate_669(G1417,G1413);
nand gate_670(G520,G1453,G1456);
not gate_671(G1457,G1453);
nand gate_672(G523,G1445,G1448);
not gate_673(G1449,G1445);
nand gate_674(G533,G1466,G1473);
nand gate_675(G536,G1458,muxed35);
nand gate_676(G496,G1418,G1425);
nand gate_677(G499,G1410,G1417);
nand gate_678(G521,G1450,G1457);
nand gate_679(G524,G1442,G1449);
nand gate_680(G534,G532,G533);
nand gate_681(G537,G535,muxed33);
nand gate_682(G497,G495,G496);
nand gate_683(G500,G498,muxed46);
nand gate_684(G522,G520,G521);
nand gate_685(G525,G523,G524);
not gate_686(G540,G534);
not gate_687(G503,G497);
not gate_688(G528,G522);
not gate_689(G669,muxed32);
buf gate_690(G672,muxed32);
not gate_691(G569,G500);
and gate_692(G588,G566,G500);
not gate_693(G618,G525);
and gate_694(G639,G615,G525);
nand gate_695(G867,G516,G564,G552,G540,G482,G528,G503,G487);
buf gate_696(G588a,G588);
buf gate_697(G588b,G588);
buf gate_698(G639a,G639);
buf gate_699(G639b,G639);
and gate_700(G675,G663,G669);
and gate_701(G688,G666,G669);
and gate_702(G696,G663,muxed31);
and gate_703(G710,G666,muxed31);
and gate_704(G73,G949,G867,G932,G932);
and gate_705(G572,G565,G569);
and gate_706(G573,G566,G569);
and gate_707(G621,G614,G618);
and gate_708(G622,G615,G618);
nand gate_709(G776,G588a,G639a,G696,G731,G958);
nand gate_710(G780,G588a,G639a,G675,G756,G958);
nand gate_711(G784,G588a,G639a,G675,G746,G958);
nand gate_712(G788,G588a,G639a,G688,G731,G958);
nand gate_713(G812,G588b,G639a,muxed30,G746,G969);
nand gate_714(G832,G588b,G639b,G696,muxed40,G969);
nand gate_715(G836,G588b,G639b,muxed30,G756,G969);
and gate_716(G1509,G588a,G639a,G696,G731,G958);
and gate_717(G1517,G588a,G639a,G675,G756,G958);
and gate_718(G1525,G588a,G639a,G675,G746,G958);
and gate_719(G1533,G588a,G639a,G688,G731,G958);
and gate_720(G1581,G588b,G639a,muxed30,G746,G969);
and gate_721(G1621,G588b,G639b,G696,muxed40,G969);
and gate_722(G1629,G588b,G639b,muxed30,G756,G969);
nand gate_723(G792,G588a,G622,G696,G756,G958);
nand gate_724(G796,G588b,G622,G696,G746,G958);
nand gate_725(G800,G588b,G622,muxed30,G731,G958);
nand gate_726(G804,G588b,G622,G675,muxed40,G958);
nand gate_727(G808,G588b,G622,G688,G756,G969);
nand gate_728(G816,G573,G639b,G696,G756,G969);
nand gate_729(G820,G573,G639b,G696,G746,G969);
nand gate_730(G824,G573,G639b,muxed30,G731,G969);
nand gate_731(G828,G573,G639b,G688,G756,G969);
nand gate_732(G871,G588b,G622,G675,G731,G979);
nand gate_733(G873,G573,G639b,G675,G731,G979);
nand gate_734(G875,G573,G622,G696,G731,G979);
nand gate_735(G877,G573,G622,G675,G756,G979);
nand gate_736(G879,G573,G622,G675,G746,G979);
nand gate_737(G881,G573,G622,G688,G731,G979);
nand gate_738(G883,G573,G621,G675,G731,G979);
nand gate_739(G885,G572,G622,G675,G731,G979);
and gate_740(G1541,G588a,G622,G696,G756,G958);
and gate_741(G1549,G588b,G622,G696,G746,G958);
and gate_742(G1557,G588b,G622,muxed30,G731,G958);
and gate_743(G1565,G588b,G622,G675,muxed40,G958);
and gate_744(G1573,G588b,G622,G688,G756,G969);
and gate_745(G1589,G573,G639b,G696,G756,G969);
and gate_746(G1597,G573,G639b,G696,G746,G969);
and gate_747(G1605,G573,G639b,muxed30,G731,G969);
and gate_748(G1613,G573,G639b,G688,G756,G969);
nand gate_749(G1,G1509,G1512);
not gate_750(G1513,G1509);
nand gate_751(G4,G1517,G1520);
not gate_752(G1521,G1517);
nand gate_753(G7,G1525,G1528);
not gate_754(G1529,G1525);
nand gate_755(G10,G1533,G1536);
not gate_756(G1537,G1533);
nand gate_757(G28,G1581,G1584);
not gate_758(G1585,G1581);
nand gate_759(G43,G1621,G1624);
not gate_760(G1625,G1621);
nand gate_761(G46,G1629,G1632);
not gate_762(G1633,G1629);
and gate_763(G886,G871,G873,G875,G877,G879,G881,G883,G885);
nand gate_764(G2,G1506,G1513);
nand gate_765(G5,G1514,G1521);
nand gate_766(G8,G1522,G1529);
nand gate_767(G11,G1530,G1537);
nand gate_768(G13,G1541,G1544);
not gate_769(G1545,G1541);
nand gate_770(G16,G1549,G1552);
not gate_771(G1553,G1549);
nand gate_772(G19,G1557,G1560);
not gate_773(G1561,G1557);
nand gate_774(G22,muxed39,G1568);
not gate_775(G1569,muxed39);
nand gate_776(G25,G1573,G1576);
not gate_777(G1577,G1573);
nand gate_778(G29,G1578,G1585);
nand gate_779(G31,G1589,muxed16);
not gate_780(G1593,G1589);
nand gate_781(G34,G1597,G1600);
not gate_782(G1601,G1597);
nand gate_783(G37,muxed29,G1608);
not gate_784(G1609,muxed29);
nand gate_785(G40,G1613,G1616);
not gate_786(G1617,G1613);
nand gate_787(G44,G1618,G1625);
nand gate_788(G47,G1626,G1633);
nand gate_789(G857,G776,G780,G784,G788,G792,muxed10,G800,G804);
nand gate_790(G860,G808,G812,G816,G820,G824,G828,G832,G836);
and gate_791(G863,G776,G780,G784,G788,G792,muxed10,G800,G804);
and gate_792(G865,G808,G812,G816,G820,G824,G828,G832,G836);
nand gate_793(G3,G1,G2);
nand gate_794(G6,G4,G5);
nand gate_795(G9,G7,muxed28);
nand gate_796(G12,G10,G11);
nand gate_797(G14,G1538,G1545);
nand gate_798(G17,G1546,G1553);
nand gate_799(G20,G1554,G1561);
nand gate_800(G23,G1562,muxed38);
nand gate_801(G26,G1570,G1577);
nand gate_802(G30,G28,G29);
nand gate_803(G32,G1586,G1593);
nand gate_804(G35,G1594,G1601);
nand gate_805(G38,G1602,muxed27);
nand gate_806(G41,G1610,G1617);
nand gate_807(G45,G43,G44);
nand gate_808(G48,G46,G47);
and gate_809(G1913,G857,G859);
and gate_810(G1921,G860,G862);
nand gate_811(G15,G13,G14);
nand gate_812(G18,G16,G17);
nand gate_813(G21,G19,G20);
nand gate_814(G24,G22,G23);
nand gate_815(G27,G25,G26);
nand gate_816(G33,G31,G32);
nand gate_817(G36,G34,G35);
nand gate_818(G39,G37,muxed4);
nand gate_819(G42,G40,G41);
and gate_820(G887,G863,G865,G886);
nand gate_821(G462,G863,G865);
and gate_822(G74,G949,G867,G952,G887);
nand gate_823(G1637,G1913,G1916);
not gate_824(G1917,G1913);
nand gate_825(G1647,G1921,G1924);
not gate_826(G1925,G1921);
nor gate_827(G75,G73,G74);
and gate_828(G1020,G457,G911,G462);
and gate_829(G1144,G469,G911,G462);
and gate_830(G1386,G475,G911,G462);
and gate_831(G1394,G478,G911,G462);
and gate_832(G1402,G459,G911,G462);
nand gate_833(G1638,G1910,G1917);
nand gate_834(G1648,G1918,G1925);
and gate_835(G1806,G472,G911,G462);
nand gate_836(G1639,G1637,G1638);
nand gate_837(G1649,G1647,G1648);
nand gate_838(G287,G1020,G1029);
nand gate_839(G350,G1144,G1153);
nand gate_840(G427,G1386,G1393);
nand gate_841(G429,G1394,G1401);
nand gate_842(G431,G1402,G1409);
not gate_843(G1028,G1020);
not gate_844(G1152,G1144);
not gate_845(G1392,G1386);
not gate_846(G1400,G1394);
not gate_847(G1408,G1402);
not gate_848(G1812,G1806);
nand gate_849(G1216,G1806,G1813);
nand gate_850(G286,G1025,G1028);
nand gate_851(G349,G1149,G1152);
nand gate_852(G426,G1389,G1392);
nand gate_853(G428,G1397,G1400);
nand gate_854(G430,G1405,G1408);
nand gate_855(G67,G1639,G1642);
not gate_856(G1643,G1639);
nand gate_857(G70,G1649,G1652);
not gate_858(G1653,G1649);
nand gate_859(G1215,G1809,G1812);
nand gate_860(G49,G286,G287);
nand gate_861(G53,G349,G350);
nand gate_862(G59,G426,G427);
nand gate_863(G61,G428,G429);
nand gate_864(G65,G430,G431);
nand gate_865(G68,G1634,G1643);
nand gate_866(G71,G1644,G1653);
nand gate_867(G1217,G1215,G1216);
and gate_868(G51,G49,G50);
and gate_869(G54,G52,G53);
and gate_870(G60,G58,G59);
and gate_871(G63,G61,G62);
and gate_872(G66,G64,G65);
nand gate_873(G69,G67,G68);
nand gate_874(G72,G70,G71);
nand gate_875(G375,G1217,G1220);
not gate_876(G1221,G1217);
nand gate_877(G376,G1212,G1221);
nand gate_878(G55,G375,muxed22);
and gate_879(G57,G55,G56);
assign muxed0 = keyinput0 ? G983 : muxed1;
assign muxed1 = keyinput1 ? G1143 : G1033;
assign muxed2 = keyinput2 ? G1139 : G296;
assign muxed3 = keyinput3 ? G1137 : G1702;
assign muxed4 = keyinput4 ? muxed26 : G1137;
assign muxed5 = keyinput5 ? G1769 : G1693;
assign muxed6 = keyinput6 ? G262 : G1202;
assign muxed7 = keyinput7 ? G261 : G1717;
assign muxed8 = keyinput8 ? G1184 : G261;
assign muxed9 = keyinput9 ? G989 : G1298;
assign muxed10 = keyinput10 ? G796 : G989;
assign muxed11 = keyinput11 ? G985 : G1216;
assign muxed12 = keyinput12 ? G990 : muxed13;
assign muxed13 = keyinput13 ? G1019 : G618;
assign muxed14 = keyinput14 ? G1015 : G988;
assign muxed15 = keyinput15 ? G1014 : G273;
assign muxed16 = keyinput16 ? G1592 : G1014;
assign muxed17 = keyinput17 ? G1685 : G1232;
assign muxed18 = keyinput18 ? G1886 : G1685;
assign muxed19 = keyinput19 ? G1681 : G1686;
assign muxed20 = keyinput20 ? G265 : G1088;
assign muxed21 = keyinput21 ? G259 : G1377;
assign muxed22 = keyinput22 ? G376 : G259;
assign muxed23 = keyinput23 ? G258 : G500;
assign muxed24 = keyinput24 ? G1050 : G258;
assign muxed25 = keyinput25 ? G1461 : muxed26;
assign muxed26 = keyinput26 ? G38 : G1700;
assign muxed27 = keyinput27 ? G1609 : G1416;
assign muxed28 = keyinput28 ? G8 : G1609;
assign muxed29 = keyinput29 ? G1605 : G1072;
assign muxed30 = keyinput30 ? G710 : G1453;
assign muxed31 = keyinput31 ? G672 : G1448;
assign muxed32 = keyinput32 ? G537 : G1332;
assign muxed33 = keyinput33 ? G536 : G231;
assign muxed34 = keyinput34 ? G549 : G536;
assign muxed35 = keyinput35 ? G1465 : G457;
assign muxed36 = keyinput36 ? G314 : G1465;
assign muxed37 = keyinput37 ? G449 : muxed38;
assign muxed38 = keyinput38 ? G1569 : G1325;
assign muxed39 = keyinput39 ? G1565 : G397;
assign muxed40 = keyinput40 ? G770 : G1693;
assign muxed41 = keyinput41 ? G722 : G433;
assign muxed42 = keyinput42 ? G561 : G639;
assign muxed43 = keyinput43 ? G560 : G1440;
assign muxed44 = keyinput44 ? G1265 : G560;
assign muxed45 = keyinput45 ? G1497 : G285;
assign muxed46 = keyinput46 ? G499 : G1497;
assign muxed47 = keyinput47 ? G1493 : G1212;
endmodule
