`timescale 1ns / 1ps
// Verilog
// c499
// Ninputs 41
// Noutputs 32
// NtotalGates 202
// XOR2 104
// AND2 40
// NOT1 40
// AND4 8
// OR4 2
// AND5 8

module top (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
                  N753,N754,N755,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
                  keyinput60, keyinput61, keyinput62, keyinput63,
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
        keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
        keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
        keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
        keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
        keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
        keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
        keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
                  keyinput144, keyinput145,
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150,
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155,
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160,
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165,
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170,
        keyinput171, keyinput172, keyinput173, keyinput174, keyinput175,
        keyinput176, keyinput177, keyinput178, keyinput179, keyinput180,
        keyinput181, keyinput182, keyinput183, keyinput184, keyinput185,
        keyinput186);

  input keyinput146, keyinput147, keyinput148, keyinput149, keyinput150;
  input keyinput151, keyinput152, keyinput153, keyinput154, keyinput155;
  input keyinput156, keyinput157, keyinput158, keyinput159, keyinput160;
  input keyinput161, keyinput162, keyinput163, keyinput164, keyinput165;
  input keyinput166, keyinput167, keyinput168, keyinput169, keyinput170;
  input keyinput171, keyinput172, keyinput173, keyinput174, keyinput175;
  input keyinput176, keyinput177, keyinput178, keyinput179, keyinput180;
  input keyinput181, keyinput182, keyinput183, keyinput184, keyinput185;
  input keyinput186;


  input keyinput64, keyinput65, keyinput66, keyinput67, keyinput68;
  input keyinput69, keyinput70, keyinput71, keyinput72, keyinput73;
  input keyinput74, keyinput75, keyinput76, keyinput77, keyinput78;
  input keyinput79, keyinput80, keyinput81, keyinput82, keyinput83;
  input keyinput84, keyinput85, keyinput86, keyinput87, keyinput88;
  input keyinput89, keyinput90, keyinput91, keyinput92, keyinput93;
  input keyinput94, keyinput95, keyinput96, keyinput97, keyinput98;
  input keyinput99, keyinput100, keyinput101, keyinput102, keyinput103;
  input keyinput104, keyinput105, keyinput106, keyinput107, keyinput108;
  input keyinput109, keyinput110, keyinput111, keyinput112, keyinput113;
  input keyinput114, keyinput115, keyinput116, keyinput117, keyinput118;
  input keyinput119, keyinput120, keyinput121, keyinput122, keyinput123;
  input keyinput124, keyinput125, keyinput126, keyinput127, keyinput128;
  input keyinput129, keyinput130, keyinput131, keyinput132, keyinput133;
  input keyinput134, keyinput135, keyinput136, keyinput137, keyinput138;
  input keyinput139, keyinput140, keyinput141, keyinput142, keyinput143;
  input keyinput144, keyinput145;

  wire KeyWire_0_1 , KeyWire_0_2;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31, keyinput32, keyinput33, keyinput34;
  input keyinput35, keyinput36, keyinput37, keyinput38, keyinput39;
  input keyinput40, keyinput41, keyinput42, keyinput43, keyinput44;
  input keyinput45, keyinput46, keyinput47, keyinput48, keyinput49;
  input keyinput50, keyinput51, keyinput52, keyinput53, keyinput54;
  input keyinput55, keyinput56, keyinput57, keyinput58, keyinput59;
  input keyinput60, keyinput61, keyinput62, keyinput63;

  wire [0:63] keyinput_Wire_0;
  wire [0:29] KeyNOTWire_0;

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;

output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723;

  xor XOR2_1 (keyinput_Wire_0[0], N1, N5);
  xor keyGate_0_0(N250, keyinput0, keyinput_Wire_0[0]);
xor XOR2_2 (N251, N9, N13);
xor XOR2_3 (N252, N17, N21);
  xor XOR2_4 (keyinput_Wire_0[1], N25, N29);
  xnor keyGate_0_1(N253, keyinput1, keyinput_Wire_0[1]);
xor XOR2_5 (N254, N33, N37);
xor XOR2_6 (N255, N41, N45);
  xor XOR2_7 (keyinput_Wire_0[2], N49, N53);
  xnor keyGate_0_2(KeyNOTWire_0[0], keyinput2, keyinput_Wire_0[2]);
  not KeyNOTGate_0_0(N256, KeyNOTWire_0[0]);
  xor XOR2_8 (keyinput_Wire_0[3], N57, N61);
  xor keyGate_0_3(KeyNOTWire_0[1], keyinput3, keyinput_Wire_0[3]);
  not KeyNOTGate_0_1(N257, KeyNOTWire_0[1]);
xor XOR2_9 (N258, N65, N69);
xor XOR2_10 (N259, N73, N77);
xor XOR2_11 (N260, N81, N85);
xor XOR2_12 (N261, N89, N93);
xor XOR2_13 (N262, N97, N101);
  xor XOR2_14 (keyinput_Wire_0[4], N105, N109);
  xor keyGate_0_4(KeyNOTWire_0[2], keyinput4, keyinput_Wire_0[4]);
  not KeyNOTGate_0_2(N263, KeyNOTWire_0[2]);
xor XOR2_15 (N264, N113, N117);
xor XOR2_16 (N265, N121, N125);
and AND2_17 (N266, N129, N137);
  and AND2_18 (keyinput_Wire_0[5], N130, N137);
  xnor keyGate_0_5(KeyNOTWire_0[3], keyinput5, keyinput_Wire_0[5]);
  not KeyNOTGate_0_3(N267, KeyNOTWire_0[3]);
and AND2_19 (N268, N131, N137);
  and AND2_20 (keyinput_Wire_0[6], N132, N137);
  xnor keyGate_0_6(N269, keyinput6, keyinput_Wire_0[6]);
and AND2_21 (N270, N133, N137);
and AND2_22 (N271, N134, N137);
and AND2_23 (N272, N135, N137);
and AND2_24 (N273, N136, N137);
xor XOR2_25 (N274, N1, N17);
  xor XOR2_26 (keyinput_Wire_0[7], N33, N49);
  xnor keyGate_0_7(N275, keyinput7, keyinput_Wire_0[7]);
xor XOR2_27 (N276, N5, N21);
  xor XOR2_28 (keyinput_Wire_0[8], N37, N53);
  xor keyGate_0_8(N277, keyinput8, keyinput_Wire_0[8]);
xor XOR2_29 (N278, N9, N25);
xor XOR2_30 (N279, N41, N57);
xor XOR2_31 (N280, N13, N29);
xor XOR2_32 (N281, N45, N61);
xor XOR2_33 (N282, N65, N81);
xor XOR2_34 (N283, N97, N113);
  xor XOR2_35 (keyinput_Wire_0[9], N69, N85);
  xnor keyGate_0_9(N284, keyinput9, keyinput_Wire_0[9]);
xor XOR2_36 (N285, N101, N117);
xor XOR2_37 (N286, N73, N89);
xor XOR2_38 (N287, N105, N121);
xor XOR2_39 (N288, N77, N93);
xor XOR2_40 (N289, N109, N125);
  xor XOR2_41 (keyinput_Wire_0[10], N250, N251);
  xnor keyGate_0_10(N290, keyinput10, keyinput_Wire_0[10]);
  xor XOR2_42 (keyinput_Wire_0[11], N252, N253);
  xor keyGate_0_11(N293, keyinput11, keyinput_Wire_0[11]);
xor XOR2_43 (N296, N254, N255);
  xor XOR2_44 (keyinput_Wire_0[12], N256, N257);
  xor keyGate_0_12(N299, keyinput12, keyinput_Wire_0[12]);
xor XOR2_45 (N302, N258, N259);
xor XOR2_46 (N305, N260, N261);
xor XOR2_47 (N308, N262, N263);
  xor XOR2_48 (keyinput_Wire_0[13], N264, N265);
  xor keyGate_0_13(KeyNOTWire_0[4], keyinput13, keyinput_Wire_0[13]);
  not KeyNOTGate_0_4(N311, KeyNOTWire_0[4]);
  xor XOR2_49 (keyinput_Wire_0[14], N274, N275);
  xnor keyGate_0_14(KeyNOTWire_0[5], keyinput14, keyinput_Wire_0[14]);
  not KeyNOTGate_0_5(N314, KeyNOTWire_0[5]);
xor XOR2_50 (N315, N276, N277);
xor XOR2_51 (N316, N278, N279);
  xor XOR2_52 (keyinput_Wire_0[15], N280, N281);
  xnor keyGate_0_15(KeyNOTWire_0[6], keyinput15, keyinput_Wire_0[15]);
  not KeyNOTGate_0_6(N317, KeyNOTWire_0[6]);
  xor XOR2_53 (keyinput_Wire_0[16], N282, N283);
  xnor keyGate_0_16(N318, keyinput16, keyinput_Wire_0[16]);
xor XOR2_54 (N319, N284, N285);
xor XOR2_55 (N320, N286, N287);
xor XOR2_56 (N321, N288, N289);
  xor XOR2_57 (keyinput_Wire_0[17], N290, N293);
  xnor keyGate_0_17(N338, keyinput17, keyinput_Wire_0[17]);
  xor XOR2_58 (keyinput_Wire_0[18], N296, N299);
  xor keyGate_0_18(N339, keyinput18, keyinput_Wire_0[18]);
  xor XOR2_59 (keyinput_Wire_0[19], N290, N296);
  xor keyGate_0_19(KeyNOTWire_0[7], keyinput19, keyinput_Wire_0[19]);
  not KeyNOTGate_0_7(N340, KeyNOTWire_0[7]);
xor XOR2_60 (N341, N293, N299);
xor XOR2_61 (N342, N302, N305);
xor XOR2_62 (N343, N308, N311);
xor XOR2_63 (N344, N302, N308);
  xor XOR2_64 (keyinput_Wire_0[20], N305, N311);
  xnor keyGate_0_20(N345, keyinput20, keyinput_Wire_0[20]);
  xor XOR2_65 (keyinput_Wire_0[21], N266, N342);
  xor keyGate_0_21(KeyNOTWire_0[8], keyinput21, keyinput_Wire_0[21]);
  not KeyNOTGate_0_8(N346, KeyNOTWire_0[8]);
xor XOR2_66 (N347, N267, N343);
xor XOR2_67 (N348, N268, N344);
xor XOR2_68 (N349, N269, N345);
xor XOR2_69 (N350, N270, N338);
xor XOR2_70 (N351, N271, N339);
xor XOR2_71 (N352, N272, N340);
xor XOR2_72 (N353, N273, N341);
  xor XOR2_73 (keyinput_Wire_0[22], N314, N346);
  xor keyGate_0_22(KeyNOTWire_0[9], keyinput22, keyinput_Wire_0[22]);
  not KeyNOTGate_0_9(N354, KeyNOTWire_0[9]);
xor XOR2_74 (N367, N315, N347);
  xor XOR2_75 (keyinput_Wire_0[23], N316, N348);
  xnor keyGate_0_23(KeyNOTWire_0[10], keyinput23, keyinput_Wire_0[23]);
  not KeyNOTGate_0_10(N380, KeyNOTWire_0[10]);
xor XOR2_76 (N393, N317, N349);
xor XOR2_77 (N406, N318, N350);
  xor XOR2_78 (keyinput_Wire_0[24], N319, N351);
  xnor keyGate_0_24(KeyNOTWire_0[11], keyinput24, keyinput_Wire_0[24]);
  not KeyNOTGate_0_11(N419, KeyNOTWire_0[11]);
xor XOR2_79 (N432, N320, N352);
xor XOR2_80 (N445, N321, N353);
not NOT1_81 (N554, N354);
not NOT1_82 (N555, N367);
not NOT1_83 (N556, N380);
not NOT1_84 (N557, N354);
not NOT1_85 (N558, N367);
not NOT1_86 (N559, N393);
  not NOT1_87 (keyinput_Wire_0[25], N354);
  xnor keyGate_0_25(N560, keyinput25, keyinput_Wire_0[25]);
  not NOT1_88 (keyinput_Wire_0[26], N380);
  xor keyGate_0_26(N561, keyinput26, keyinput_Wire_0[26]);
  not NOT1_89 (keyinput_Wire_0[27], N393);
  xnor keyGate_0_27(N562, keyinput27, keyinput_Wire_0[27]);
not NOT1_90 (N563, N367);
not NOT1_91 (N564, N380);
not NOT1_92 (N565, N393);
not NOT1_93 (N566, N419);
  not NOT1_94 (keyinput_Wire_0[28], N445);
  xor keyGate_0_28(KeyNOTWire_0[12], keyinput28, keyinput_Wire_0[28]);
  not KeyNOTGate_0_12(N567, KeyNOTWire_0[12]);
not NOT1_95 (N568, N419);
not NOT1_96 (N569, N432);
not NOT1_97 (N570, N406);
  not NOT1_98 (keyinput_Wire_0[29], N445);
  xnor keyGate_0_29(KeyNOTWire_0[13], keyinput29, keyinput_Wire_0[29]);
  not KeyNOTGate_0_13(N571, KeyNOTWire_0[13]);
not NOT1_99 (N572, N406);
not NOT1_100 (N573, N432);
not NOT1_101 (N574, N406);
not NOT1_102 (N575, N419);
  not NOT1_103 (keyinput_Wire_0[30], N432);
  xor keyGate_0_30(N576, keyinput30, keyinput_Wire_0[30]);
not NOT1_104 (N577, N406);
  not NOT1_105 (keyinput_Wire_0[31], N419);
  xor keyGate_0_31(N578, keyinput31, keyinput_Wire_0[31]);
not NOT1_106 (N579, N445);
not NOT1_107 (N580, N406);
  not NOT1_108 (keyinput_Wire_0[32], N432);
  xor keyGate_0_32(N581, keyinput32, keyinput_Wire_0[32]);
  not NOT1_109 (keyinput_Wire_0[33], N445);
  xnor keyGate_0_33(KeyNOTWire_0[14], keyinput33, keyinput_Wire_0[33]);
  not KeyNOTGate_0_14(N582, KeyNOTWire_0[14]);
  not NOT1_110 (keyinput_Wire_0[34], N419);
  xor keyGate_0_34(N583, keyinput34, keyinput_Wire_0[34]);
not NOT1_111 (N584, N432);
not NOT1_112 (N585, N445);
  not NOT1_113 (keyinput_Wire_0[35], N367);
  xor keyGate_0_35(KeyNOTWire_0[15], keyinput35, keyinput_Wire_0[35]);
  not KeyNOTGate_0_15(N586, KeyNOTWire_0[15]);
not NOT1_114 (N587, N393);
not NOT1_115 (N588, N367);
  not NOT1_116 (keyinput_Wire_0[36], N380);
  xor keyGate_0_36(KeyNOTWire_0[16], keyinput36, keyinput_Wire_0[36]);
  not KeyNOTGate_0_16(N589, KeyNOTWire_0[16]);
not NOT1_117 (N590, N354);
not NOT1_118 (N591, N393);
not NOT1_119 (N592, N354);
not NOT1_120 (N593, N380);
  and AND4_121 (keyinput_Wire_0[37], N554, N555, N556, N393);
  xnor keyGate_0_37(KeyNOTWire_0[17], keyinput37, keyinput_Wire_0[37]);
  not KeyNOTGate_0_17(N594, KeyNOTWire_0[17]);
and AND4_122 (N595, N557, N558, N380, N559);
and AND4_123 (N596, N560, N367, N561, N562);
and AND4_124 (N597, N354, N563, N564, N565);
  and AND4_125 (keyinput_Wire_0[38], N574, N575, N576, N445);
  xor keyGate_0_38(N598, keyinput38, keyinput_Wire_0[38]);
and AND4_126 (N599, N577, N578, N432, N579);
  and AND4_127 (keyinput_Wire_0[39], N580, N419, N581, N582);
  xnor keyGate_0_39(N600, keyinput39, keyinput_Wire_0[39]);
and AND4_128 (N601, N406, N583, N584, N585);
or OR4_129 (N602, N594, N595, N596, N597);
  or OR4_130 (keyinput_Wire_0[40], N598, N599, N600, N601);
  xor keyGate_0_40(N607, keyinput40, keyinput_Wire_0[40]);
and AND5_131 (N620, N406, N566, N432, N567, N602);
and AND5_132 (N625, N406, N568, N569, N445, N602);
and AND5_133 (N630, N570, N419, N432, N571, N602);
and AND5_134 (N635, N572, N419, N573, N445, N602);
and AND5_135 (N640, N354, N586, N380, N587, N607);
and AND5_136 (N645, N354, N588, N589, N393, N607);
  and AND5_137 (keyinput_Wire_0[41], N590, N367, N380, N591, N607);
  xor keyGate_0_41(KeyNOTWire_0[18], keyinput41, keyinput_Wire_0[41]);
  not KeyNOTGate_0_18(N650, KeyNOTWire_0[18]);
and AND5_138 (N655, N592, N367, N593, N393, N607);
and AND2_139 (N692, N354, N620);
and AND2_140 (N693, N367, N620);
  and AND2_141 (keyinput_Wire_0[42], N380, N620);
  xor keyGate_0_42(KeyNOTWire_0[19], keyinput42, keyinput_Wire_0[42]);
  not KeyNOTGate_0_19(N694, KeyNOTWire_0[19]);
and AND2_142 (N695, N393, N620);
  and AND2_143 (keyinput_Wire_0[43], N354, N625);
  xnor keyGate_0_43(N696, keyinput43, keyinput_Wire_0[43]);
and AND2_144 (N697, N367, N625);
  and AND2_145 (keyinput_Wire_0[44], N380, N625);
  xor keyGate_0_44(KeyNOTWire_0[20], keyinput44, keyinput_Wire_0[44]);
  not KeyNOTGate_0_20(N698, KeyNOTWire_0[20]);
  and AND2_146 (keyinput_Wire_0[45], N393, N625);
  xor keyGate_0_45(KeyNOTWire_0[21], keyinput45, keyinput_Wire_0[45]);
  not KeyNOTGate_0_21(N699, KeyNOTWire_0[21]);
and AND2_147 (N700, N354, N630);
  and AND2_148 (keyinput_Wire_0[46], N367, N630);
  xnor keyGate_0_46(N701, keyinput46, keyinput_Wire_0[46]);
  and AND2_149 (keyinput_Wire_0[47], N380, N630);
  xnor keyGate_0_47(N702, keyinput47, keyinput_Wire_0[47]);
and AND2_150 (N703, N393, N630);
and AND2_151 (N704, N354, N635);
  and AND2_152 (keyinput_Wire_0[48], N367, N635);
  xor keyGate_0_48(KeyNOTWire_0[22], keyinput48, keyinput_Wire_0[48]);
  not KeyNOTGate_0_22(N705, KeyNOTWire_0[22]);
  and AND2_153 (keyinput_Wire_0[49], N380, N635);
  xnor keyGate_0_49(KeyNOTWire_0[23], keyinput49, keyinput_Wire_0[49]);
  not KeyNOTGate_0_23(N706, KeyNOTWire_0[23]);
and AND2_154 (N707, N393, N635);
and AND2_155 (N708, N406, N640);
and AND2_156 (N709, N419, N640);
  and AND2_157 (keyinput_Wire_0[50], N432, N640);
  xnor keyGate_0_50(KeyNOTWire_0[24], keyinput50, keyinput_Wire_0[50]);
  not KeyNOTGate_0_24(N710, KeyNOTWire_0[24]);
  and AND2_158 (keyinput_Wire_0[51], N445, N640);
  xnor keyGate_0_51(KeyNOTWire_0[25], keyinput51, keyinput_Wire_0[51]);
  not KeyNOTGate_0_25(N711, KeyNOTWire_0[25]);
and AND2_159 (N712, N406, N645);
and AND2_160 (N713, N419, N645);
and AND2_161 (N714, N432, N645);
and AND2_162 (N715, N445, N645);
and AND2_163 (N716, N406, N650);
and AND2_164 (N717, N419, N650);
and AND2_165 (N718, N432, N650);
and AND2_166 (N719, N445, N650);
  and AND2_167 (keyinput_Wire_0[52], N406, N655);
  xnor keyGate_0_52(N720, keyinput52, keyinput_Wire_0[52]);
and AND2_168 (N721, N419, N655);
and AND2_169 (N722, N432, N655);
and AND2_170 (N723, N445, N655);
  xor XOR2_171 (keyinput_Wire_0[53], N1, N692);
  xnor keyGate_0_53(KeyNOTWire_0[26], keyinput53, keyinput_Wire_0[53]);
  not KeyNOTGate_0_26(N724, KeyNOTWire_0[26]);
xor XOR2_172 (N725, N5, N693);
xor XOR2_173 (N726, N9, N694);
xor XOR2_174 (N727, N13, N695);
  xor XOR2_175 (keyinput_Wire_0[54], N17, N696);
  xor keyGate_0_54(KeyNOTWire_0[27], keyinput54, keyinput_Wire_0[54]);
  not KeyNOTGate_0_27(N728, KeyNOTWire_0[27]);
xor XOR2_176 (N729, N21, N697);
  xor XOR2_177 (keyinput_Wire_0[55], N25, N698);
  xor keyGate_0_55(N730, keyinput55, keyinput_Wire_0[55]);
xor XOR2_178 (N731, N29, N699);
xor XOR2_179 (N732, N33, N700);
xor XOR2_180 (N733, N37, N701);
xor XOR2_181 (N734, N41, N702);
  xor XOR2_182 (keyinput_Wire_0[56], N45, N703);
  xor keyGate_0_56(N735, keyinput56, keyinput_Wire_0[56]);
xor XOR2_183 (N736, N49, N704);
xor XOR2_184 (N737, N53, N705);
  xor XOR2_185 (keyinput_Wire_0[57], N57, N706);
  xor keyGate_0_57(N738, keyinput57, keyinput_Wire_0[57]);
xor XOR2_186 (KeyWire_0_1, N61, N707);
  xor flip_it (N739, KeyWire_0_1, KeyWire_0_2 );
xor XOR2_187 (N740, N65, N708);
  xor XOR2_188 (keyinput_Wire_0[58], N69, N709);
  xor keyGate_0_58(KeyNOTWire_0[28], keyinput58, keyinput_Wire_0[58]);
  not KeyNOTGate_0_28(N741, KeyNOTWire_0[28]);
xor XOR2_189 (N742, N73, N710);
  xor XOR2_190 (keyinput_Wire_0[59], N77, N711);
  xnor keyGate_0_59(N743, keyinput59, keyinput_Wire_0[59]);
  xor XOR2_191 (keyinput_Wire_0[60], N81, N712);
  xnor keyGate_0_60(N744, keyinput60, keyinput_Wire_0[60]);
  xor XOR2_192 (keyinput_Wire_0[61], N85, N713);
  xor keyGate_0_61(N745, keyinput61, keyinput_Wire_0[61]);
  xor XOR2_193 (keyinput_Wire_0[62], N89, N714);
  xnor keyGate_0_62(KeyNOTWire_0[29], keyinput62, keyinput_Wire_0[62]);
  not KeyNOTGate_0_29(N746, KeyNOTWire_0[29]);
xor XOR2_194 (N747, N93, N715);
xor XOR2_195 (N748, N97, N716);
  xor XOR2_196 (keyinput_Wire_0[63], N101, N717);
  xnor keyGate_0_63(N749, keyinput63, keyinput_Wire_0[63]);
xor XOR2_197 (N750, N105, N718);
xor XOR2_198 (N751, N109, N719);
xor XOR2_199 (N752, N113, N720);
xor XOR2_200 (N753, N117, N721);
xor XOR2_201 (N754, N121, N722);
xor XOR2_202 (N755, N125, N723);

AntiSAT some_name( KeyWire_0_2, N136, N121, N113, N137, N129, N33, N41, N125, N9, N117, N85, N37, N132, N73, N135, N1, N81, N77, N45, N105, N93, N61, N5, N13, N131, N21, N57, N133, N109, N134, N65, N101, N89, N97, N49, N29, N53, N25, N17, N130, N69, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145,
       keyinput146, keyinput147, keyinput148, keyinput149, keyinput150,
       keyinput151, keyinput152, keyinput153, keyinput154, keyinput155,
       keyinput156, keyinput157, keyinput158, keyinput159, keyinput160,
       keyinput161, keyinput162, keyinput163, keyinput164, keyinput165,
       keyinput166, keyinput167, keyinput168, keyinput169, keyinput170,
       keyinput171, keyinput172, keyinput173, keyinput174, keyinput175,
       keyinput176, keyinput177, keyinput178, keyinput179, keyinput180,
       keyinput181, keyinput182, keyinput183, keyinput184, keyinput185,
       keyinput186);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N136, N121, N113, N137, N129, N33, N41, N125, N9, N117, N85, N37, N132, N73, N135, N1, N81, N77, N45, N105, N93, N61, N5, N13, N131, N21, N57, N133, N109, N134, N65, N101, N89, N97, N49, N29, N53, N25, N17, N130, N69, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145 ,
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150,
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155,
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160,
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165,
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170,
        keyinput171, keyinput172, keyinput173, keyinput174, keyinput175,
        keyinput176, keyinput177, keyinput178, keyinput179, keyinput180,
        keyinput181, keyinput182, keyinput183, keyinput184, keyinput185,
        keyinput186);

  input keyinput146, keyinput147, keyinput148, keyinput149, keyinput150;
  input keyinput151, keyinput152, keyinput153, keyinput154, keyinput155;
  input keyinput156, keyinput157, keyinput158, keyinput159, keyinput160;
  input keyinput161, keyinput162, keyinput163, keyinput164, keyinput165;
  input keyinput166, keyinput167, keyinput168, keyinput169, keyinput170;
  input keyinput171, keyinput172, keyinput173, keyinput174, keyinput175;
  input keyinput176, keyinput177, keyinput178, keyinput179, keyinput180;
  input keyinput181, keyinput182, keyinput183, keyinput184, keyinput185;
  input keyinput186;

  wire [0:40] keyNTin_Wire_1;
  wire [0:14] KeyNOTWire_1;

  input N136, N121, N113, N137, N129, N33, N41, N125, N9, N117, N85, N37, N132, N73, N135, N1, N81, N77, N45, N105, N93, N61, N5, N13, N131, N21, N57, N133, N109, N134, N65, N101, N89, N97, N49, N29, N53, N25, N17, N130, N69;
  input keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83 ;

  xnor KeyGate0 (newWire_0, N136, keyinput64);
  xor  KeyGate1 (newWire_1, N121, keyinput65);
  xnor KeyGate2 (keyNTin_Wire_1[0], N113, keyinput66);
  xnor keyNTinGate_1_0(newWire_2, keyinput146, keyNTin_Wire_1[0]);
  xor  KeyGate3 (keyNTin_Wire_1[1], N137, keyinput67);
  xnor keyNTinGate_1_1(newWire_3, keyinput147, keyNTin_Wire_1[1]);
  xnor KeyGate4 (keyNTin_Wire_1[2], N129, keyinput68);
  xor keyNTinGate_1_2(newWire_4, keyinput148, keyNTin_Wire_1[2]);
  xor  KeyGate5 (newWire_5, N33, keyinput69);
  xnor KeyGate6 (newWire_6, N41, keyinput70);
  xor  KeyGate7 (newWire_7, N125, keyinput71);
  xor  KeyGate8 (keyNTin_Wire_1[3], N9, keyinput72);
  xnor keyNTinGate_1_3(newWire_8, keyinput149, keyNTin_Wire_1[3]);
  xor  KeyGate9 (keyNTin_Wire_1[4], N117, keyinput73);
  xnor keyNTinGate_1_4(newWire_9, keyinput150, keyNTin_Wire_1[4]);
  xnor KeyGate10 (newWire_10, N85, keyinput74);
  xor  KeyGate11 (keyNTin_Wire_1[5], N37, keyinput75);
  xnor keyNTinGate_1_5(KeyNOTWire_1[0], keyinput151, keyNTin_Wire_1[5]);
  not KeyNOTGate_1_0(newWire_11, KeyNOTWire_1[0]);
  xor  KeyGate12 (keyNTin_Wire_1[6], N132, keyinput76);
  xnor keyNTinGate_1_6(newWire_12, keyinput152, keyNTin_Wire_1[6]);
  xor  KeyGate13 (newWire_13, N73, keyinput77);
  xor  KeyGate14 (newWire_14, N135, keyinput78);
  xor  KeyGate15 (newWire_15, N1, keyinput79);
  xor  KeyGate16 (newWire_16, N81, keyinput80);
  xor  KeyGate17 (keyNTin_Wire_1[7], N77, keyinput81);
  xnor keyNTinGate_1_7(newWire_17, keyinput153, keyNTin_Wire_1[7]);
  xor  KeyGate18 (newWire_18, N45, keyinput82);
  xor  KeyGate19 (keyNTin_Wire_1[8], N105, keyinput83);
  xnor keyNTinGate_1_8(KeyNOTWire_1[1], keyinput154, keyNTin_Wire_1[8]);
  not KeyNOTGate_1_1(newWire_19, KeyNOTWire_1[1]);
  xor  KeyGate20 (keyNTin_Wire_1[9], N93, keyinput84);
  xor keyNTinGate_1_9(newWire_20, keyinput155, keyNTin_Wire_1[9]);
  xor  KeyGate21 (newWire_21, N61, keyinput85);
  xnor KeyGate22 (keyNTin_Wire_1[10], N5, keyinput86);
  xnor keyNTinGate_1_10(KeyNOTWire_1[2], keyinput156, keyNTin_Wire_1[10]);
  not KeyNOTGate_1_2(newWire_22, KeyNOTWire_1[2]);
  xnor KeyGate23 (newWire_23, N13, keyinput87);
  xnor KeyGate24 (keyNTin_Wire_1[11], N131, keyinput88);
  xnor keyNTinGate_1_11(KeyNOTWire_1[3], keyinput157, keyNTin_Wire_1[11]);
  not KeyNOTGate_1_3(newWire_24, KeyNOTWire_1[3]);
  xnor KeyGate25 (newWire_25, N21, keyinput89);
  xnor KeyGate26 (newWire_26, N57, keyinput90);
  xor  KeyGate27 (newWire_27, N133, keyinput91);
  xnor KeyGate28 (newWire_28, N109, keyinput92);
  xor  KeyGate29 (newWire_29, N134, keyinput93);
  xor  KeyGate30 (newWire_30, N65, keyinput94);
  xor  KeyGate31 (keyNTin_Wire_1[12], N101, keyinput95);
  xor keyNTinGate_1_12(newWire_31, keyinput158, keyNTin_Wire_1[12]);
  xnor KeyGate32 (newWire_32, N89, keyinput96);
  xor  KeyGate33 (keyNTin_Wire_1[13], N97, keyinput97);
  xor keyNTinGate_1_13(newWire_33, keyinput159, keyNTin_Wire_1[13]);
  xor  KeyGate34 (keyNTin_Wire_1[14], N49, keyinput98);
  xnor keyNTinGate_1_14(newWire_34, keyinput160, keyNTin_Wire_1[14]);
  xor  KeyGate35 (keyNTin_Wire_1[15], N29, keyinput99);
  xor keyNTinGate_1_15(newWire_35, keyinput161, keyNTin_Wire_1[15]);
  xnor KeyGate36 (keyNTin_Wire_1[16], N53, keyinput100);
  xor keyNTinGate_1_16(newWire_36, keyinput162, keyNTin_Wire_1[16]);
  xor  KeyGate37 (newWire_37, N25, keyinput101);
  xnor KeyGate38 (newWire_38, N17, keyinput102);
  xnor KeyGate39 (keyNTin_Wire_1[17], N130, keyinput103);
  xor keyNTinGate_1_17(newWire_39, keyinput163, keyNTin_Wire_1[17]);
  xor  KeyGate40 (keyNTin_Wire_1[18], N69, keyinput104);
  xor keyNTinGate_1_18(newWire_40, keyinput164, keyNTin_Wire_1[18]);
  xor  KeyGate41 (keyNTin_Wire_1[19], N136, keyinput105);
  xnor keyNTinGate_1_19(KeyNOTWire_1[4], keyinput165, keyNTin_Wire_1[19]);
  not KeyNOTGate_1_4(newWire_41, KeyNOTWire_1[4]);
  xor  KeyGate42 (newWire_42, N121, keyinput106);
  xor  KeyGate43 (newWire_43, N113, keyinput107);
  xnor KeyGate44 (keyNTin_Wire_1[20], N137, keyinput108);
  xor keyNTinGate_1_20(newWire_44, keyinput166, keyNTin_Wire_1[20]);
  xor  KeyGate45 (newWire_45, N129, keyinput109);
  xor  KeyGate46 (newWire_46, N33, keyinput110);
  xor  KeyGate47 (newWire_47, N41, keyinput111);
  xnor KeyGate48 (newWire_48, N125, keyinput112);
  xnor KeyGate49 (keyNTin_Wire_1[21], N9, keyinput113);
  xnor keyNTinGate_1_21(KeyNOTWire_1[5], keyinput167, keyNTin_Wire_1[21]);
  not KeyNOTGate_1_5(newWire_49, KeyNOTWire_1[5]);
  xor  KeyGate50 (newWire_50, N117, keyinput114);
  xor  KeyGate51 (newWire_51, N85, keyinput115);
  xnor KeyGate52 (keyNTin_Wire_1[22], N37, keyinput116);
  xnor keyNTinGate_1_22(newWire_52, keyinput168, keyNTin_Wire_1[22]);
  xnor KeyGate53 (keyNTin_Wire_1[23], N132, keyinput117);
  xnor keyNTinGate_1_23(KeyNOTWire_1[6], keyinput169, keyNTin_Wire_1[23]);
  not KeyNOTGate_1_6(newWire_53, KeyNOTWire_1[6]);
  xnor KeyGate54 (keyNTin_Wire_1[24], N73, keyinput118);
  xor keyNTinGate_1_24(newWire_54, keyinput170, keyNTin_Wire_1[24]);
  xnor KeyGate55 (keyNTin_Wire_1[25], N135, keyinput119);
  xnor keyNTinGate_1_25(KeyNOTWire_1[7], keyinput171, keyNTin_Wire_1[25]);
  not KeyNOTGate_1_7(newWire_55, KeyNOTWire_1[7]);
  xnor KeyGate56 (keyNTin_Wire_1[26], N1, keyinput120);
  xor keyNTinGate_1_26(KeyNOTWire_1[8], keyinput172, keyNTin_Wire_1[26]);
  not KeyNOTGate_1_8(newWire_56, KeyNOTWire_1[8]);
  xnor KeyGate57 (newWire_57, N81, keyinput121);
  xor  KeyGate58 (newWire_58, N77, keyinput122);
  xor  KeyGate59 (newWire_59, N45, keyinput123);
  xor  KeyGate60 (newWire_60, N105, keyinput124);
  xor  KeyGate61 (keyNTin_Wire_1[27], N93, keyinput125);
  xnor keyNTinGate_1_27(KeyNOTWire_1[9], keyinput173, keyNTin_Wire_1[27]);
  not KeyNOTGate_1_9(newWire_61, KeyNOTWire_1[9]);
  xnor KeyGate62 (keyNTin_Wire_1[28], N61, keyinput126);
  xor keyNTinGate_1_28(newWire_62, keyinput174, keyNTin_Wire_1[28]);
  xnor KeyGate63 (keyNTin_Wire_1[29], N5, keyinput127);
  xor keyNTinGate_1_29(newWire_63, keyinput175, keyNTin_Wire_1[29]);
  xor  KeyGate64 (newWire_64, N13, keyinput128);
  xor  KeyGate65 (keyNTin_Wire_1[30], N131, keyinput129);
  xor keyNTinGate_1_30(KeyNOTWire_1[10], keyinput176, keyNTin_Wire_1[30]);
  not KeyNOTGate_1_10(newWire_65, KeyNOTWire_1[10]);
  xor  KeyGate66 (keyNTin_Wire_1[31], N21, keyinput130);
  xor keyNTinGate_1_31(KeyNOTWire_1[11], keyinput177, keyNTin_Wire_1[31]);
  not KeyNOTGate_1_11(newWire_66, KeyNOTWire_1[11]);
  xnor KeyGate67 (newWire_67, N57, keyinput131);
  xnor KeyGate68 (newWire_68, N133, keyinput132);
  xnor KeyGate69 (keyNTin_Wire_1[32], N109, keyinput133);
  xor keyNTinGate_1_32(newWire_69, keyinput178, keyNTin_Wire_1[32]);
  xor  KeyGate70 (keyNTin_Wire_1[33], N134, keyinput134);
  xnor keyNTinGate_1_33(newWire_70, keyinput179, keyNTin_Wire_1[33]);
  xor  KeyGate71 (keyNTin_Wire_1[34], N65, keyinput135);
  xnor keyNTinGate_1_34(newWire_71, keyinput180, keyNTin_Wire_1[34]);
  xor  KeyGate72 (newWire_72, N101, keyinput136);
  xnor KeyGate73 (newWire_73, N89, keyinput137);
  xnor KeyGate74 (newWire_74, N97, keyinput138);
  xor  KeyGate75 (newWire_75, N49, keyinput139);
  xnor KeyGate76 (keyNTin_Wire_1[35], N29, keyinput140);
  xnor keyNTinGate_1_35(KeyNOTWire_1[12], keyinput181, keyNTin_Wire_1[35]);
  not KeyNOTGate_1_12(newWire_76, KeyNOTWire_1[12]);
  xor  KeyGate77 (keyNTin_Wire_1[36], N53, keyinput141);
  xnor keyNTinGate_1_36(newWire_77, keyinput182, keyNTin_Wire_1[36]);
  xor  KeyGate78 (newWire_78, N25, keyinput142);
  xor  KeyGate79 (keyNTin_Wire_1[37], N17, keyinput143);
  xor keyNTinGate_1_37(newWire_79, keyinput183, keyNTin_Wire_1[37]);
  xnor KeyGate80 (newWire_80, N130, keyinput144);
  xnor KeyGate81 (keyNTin_Wire_1[38], N69, keyinput145);
  xnor keyNTinGate_1_38(KeyNOTWire_1[13], keyinput184, keyNTin_Wire_1[38]);
  not KeyNOTGate_1_13(newWire_81, KeyNOTWire_1[13]);
  and some_function (keyNTin_Wire_1[39], newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40 );
  xnor keyNTinGate_1_39(newWire_82, keyinput185, keyNTin_Wire_1[39]);
  nand compl_function (keyNTin_Wire_1[40], newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81);
  xor keyNTinGate_1_40(KeyNOTWire_1[14], keyinput186, keyNTin_Wire_1[40]);
  not KeyNOTGate_1_14(newWire_83, KeyNOTWire_1[14]);
  and finalAND (KeyWire_0_2, newWire_82, newWire_83);

endmodule /* AntiSAT */
