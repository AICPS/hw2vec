// Verilog File 
module top (Gid0,Gid1,Gid2,Gid3,Gid4,Gid5,Gid6,Gid7,Gid8,
Gid9,Gid10,Gid11,Gid12,Gid13,Gid14,Gid15,Gid16,Gid17,Gid18,
Gid19,Gid20,Gid21,Gid22,Gid23,Gid24,Gid25,Gid26,Gid27,Gid28,
Gid29,Gid30,Gid31,Gic0,Gic1,Gic2,Gic3,Gic4,Gic5,Gic6,
Gic7,Gr,God0,God1,God2,God3,God4,God5,God6,God7,
God8,God9,God10,God11,God12,God13,God14,God15,God16,God17,
God18,God19,God20,God21,God22,God23,God24,God25,God26,God27,
God28,God29,God30,God31,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,
keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,
keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,
keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,keyinput35,
keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,keyinput45,
keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,keyinput55,
keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,keyinput65,
keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,keyinput75,
keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,keyinput85,
keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,keyinput95,
keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103);

input Gid0,Gid1,Gid2,Gid3,Gid4,Gid5,Gid6,Gid7,Gid8,
Gid9,Gid10,Gid11,Gid12,Gid13,Gid14,Gid15,Gid16,Gid17,Gid18,
Gid19,Gid20,Gid21,Gid22,Gid23,Gid24,Gid25,Gid26,Gid27,Gid28,
Gid29,Gid30,Gid31,Gic0,Gic1,Gic2,Gic3,Gic4,Gic5,Gic6,
Gic7,Gr,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,
keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,
keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,
keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,
keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,
keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,keyinput55,keyinput56,keyinput57,
keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,keyinput65,keyinput66,keyinput67,
keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,keyinput75,keyinput76,keyinput77,
keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,keyinput85,keyinput86,keyinput87,
keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,keyinput95,keyinput96,keyinput97,
keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103;

output God0,God1,God2,God3,God4,God5,God6,God7,God8,
God9,God10,God11,God12,God13,God14,God15,God16,God17,God18,
God19,God20,God21,God22,God23,God24,God25,God26,God27,God28,
God29,God30,God31;

wire Gxa0,Gxa1,Gxa2,Gxa3,Gxa4,Gxa5,Gxa6,Gxa7,Gxa8,
Gxa9,Gxa10,Gxa11,Gxa12,Gxa13,Gxa14,Gxa15,Gh0,Gh1,Gh2,
Gh3,Gh4,Gh5,Gh6,Gh7,Gxb0,Gxc0,Gxb1,Gxc1,Gxb2,
Gxc2,Gxb3,Gxc3,Gxb4,Gxc4,Gxb5,Gxc5,Gxb6,Gxc6,Gxb7,
Gxc7,Gf0,Gf1,Gf2,Gf3,Gf4,Gf5,Gf6,Gf7,Gxe0,
Gxe1,Gxe2,Gxe3,Gxe4,Gxe5,Gxe6,Gxe7,Gg0,Gg1,Gg2,
Gg3,Gg4,Gg5,Gg6,Gg7,Gxd0,Gxd1,Gxd2,Gxd3,Gxd4,
Gxd5,Gxd6,Gxd7,Gs0,Gs1,Gs2,Gs3,Gs4,Gs5,Gs6,
Gs7,Gy0a,Gy1a,Gy2a,Gy0b,Gy1b,Gy3b,Gy0c,Gy2c,Gy3c,
Gy1d,Gy2d,Gy3d,Gy5i,Gy7i,Gy5j,Gy6j,Gy4k,Gy7k,Gy4l,
Gy6l,Gy4a,Gy5a,Gy6a,Gy4b,Gy5b,Gy7b,Gy4c,Gy6c,Gy7c,
Gy5d,Gy6d,Gy7d,Gy1i,Gy3i,Gy1j,Gy2j,Gy0k,Gy3k,Gy0l,
Gy2l,Gt0,Gt1,Gt2,Gt3,Gt4,Gt5,Gt6,Gt7,Gu0,
Gu1,Gwa,Gwb,Gwc,Gwd,Gwe,Gwf,Gwg,Gwh,Ge0,
Ge1,Ge2,Ge3,Ge4,Ge5,Ge6,Ge7,Ge8,Ge9,Ge10,
Ge11,Ge12,Ge13,Ge14,Ge15,Ge16,Ge17,Ge18,Ge19,Ge20,
Ge21,Ge22,Ge23,Ge24,Ge25,Ge26,Ge27,Ge28,Ge29,Ge30,
Ge31,muxed0,muxed1,muxed2,muxed3,muxed4,muxed5,muxed6,muxed7,muxed8,
muxed9,muxed10,muxed11,muxed12,muxed13,muxed14,muxed15,muxed16,muxed17,muxed18,
muxed19,muxed20,muxed21,muxed22,muxed23,muxed24,muxed25,muxed26,muxed27,muxed28,
muxed29,muxed30,muxed31,muxed32,muxed33,muxed34,muxed35,muxed36,muxed37,muxed38,
muxed39,muxed40,muxed41,muxed42,muxed43,muxed44,muxed45,muxed46,muxed47,muxed48,
muxed49,muxed50,muxed51,muxed52,muxed53,muxed54,muxed55,muxed56,muxed57,muxed58,
muxed59,muxed60,muxed61,muxed62,muxed63,muxed64,muxed65,muxed66,muxed67,muxed68,
muxed69,muxed70,muxed71,muxed72,muxed73,muxed74,muxed75,muxed76,muxed77,muxed78,
muxed79,muxed80,muxed81,muxed82,muxed83,muxed84,muxed85,muxed86,muxed87,muxed88,
muxed89,muxed90,muxed91,muxed92,muxed93,muxed94,muxed95,muxed96,muxed97,muxed98,
muxed99,muxed100,muxed101,muxed102,muxed103;
xor gate_0(Gxa0,Gid0,Gid1);
xor gate_1(Gxa1,Gid2,Gid3);
xor gate_2(Gxa2,Gid4,Gid5);
xor gate_3(Gxa3,Gid6,Gid7);
xor gate_4(Gxa4,Gid8,Gid9);
xor gate_5(Gxa5,Gid10,Gid11);
xor gate_6(Gxa6,Gid12,Gid13);
xor gate_7(Gxa7,Gid14,Gid15);
xor gate_8(Gxa8,Gid16,Gid17);
xor gate_9(Gxa9,Gid18,Gid19);
xor gate_10(Gxa10,Gid20,Gid21);
xor gate_11(Gxa11,Gid22,Gid23);
xor gate_12(Gxa12,muxed53,Gid25);
xor gate_13(Gxa13,Gid26,Gid27);
xor gate_14(Gxa14,Gid28,Gid29);
xor gate_15(Gxa15,Gid30,Gid31);
and gate_16(Gh0,muxed41,Gr);
and gate_17(Gh1,Gic1,Gr);
and gate_18(Gh2,Gic2,Gr);
and gate_19(Gh3,Gic3,Gr);
and gate_20(Gh4,muxed0,Gr);
and gate_21(Gh5,Gic5,Gr);
and gate_22(Gh6,Gic6,Gr);
and gate_23(Gh7,Gic7,Gr);
xor gate_24(Gxb0,Gid0,Gid4);
xor gate_25(Gxc0,Gid8,Gid12);
xor gate_26(Gxb1,Gid1,Gid5);
xor gate_27(Gxc1,Gid9,Gid13);
xor gate_28(Gxb2,Gid2,Gid6);
xor gate_29(Gxc2,Gid10,Gid14);
xor gate_30(Gxb3,Gid3,Gid7);
xor gate_31(Gxc3,Gid11,Gid15);
xor gate_32(Gxb4,Gid16,Gid20);
xor gate_33(Gxc4,muxed53,Gid28);
xor gate_34(Gxb5,Gid17,Gid21);
xor gate_35(Gxc5,Gid25,Gid29);
xor gate_36(Gxb6,Gid18,Gid22);
xor gate_37(Gxc6,Gid26,Gid30);
xor gate_38(Gxb7,Gid19,Gid23);
xor gate_39(Gxc7,Gid27,Gid31);
xor gate_40(Gf0,muxed75,Gxa1);
xor gate_41(Gf1,Gxa2,Gxa3);
xor gate_42(Gf2,Gxa4,muxed54);
xor gate_43(Gf3,Gxa6,Gxa7);
xor gate_44(Gf4,Gxa8,muxed92);
xor gate_45(Gf5,Gxa10,Gxa11);
xor gate_46(Gf6,muxed62,Gxa13);
xor gate_47(Gf7,muxed13,Gxa15);
xor gate_48(Gxe0,Gxb0,Gxc0);
xor gate_49(Gxe1,Gxb1,Gxc1);
xor gate_50(Gxe2,Gxb2,Gxc2);
xor gate_51(Gxe3,Gxb3,Gxc3);
xor gate_52(Gxe4,Gxb4,Gxc4);
xor gate_53(Gxe5,Gxb5,Gxc5);
xor gate_54(Gxe6,Gxb6,Gxc6);
xor gate_55(Gxe7,Gxb7,Gxc7);
xor gate_56(Gg0,muxed74,Gf1);
xor gate_57(Gg1,Gf2,Gf3);
xor gate_58(Gg2,muxed74,Gf2);
xor gate_59(Gg3,Gf1,Gf3);
xor gate_60(Gg4,Gf4,Gf5);
xor gate_61(Gg5,muxed86,Gf7);
xor gate_62(Gg6,Gf4,muxed86);
xor gate_63(Gg7,Gf5,Gf7);
xor gate_64(Gxd0,muxed51,Gg4);
xor gate_65(Gxd1,Gh1,Gg5);
xor gate_66(Gxd2,Gh2,muxed34);
xor gate_67(Gxd3,Gh3,Gg7);
xor gate_68(Gxd4,muxed80,Gg0);
xor gate_69(Gxd5,muxed103,Gg1);
xor gate_70(Gxd6,Gh6,muxed72);
xor gate_71(Gxd7,Gh7,Gg3);
xor gate_72(Gs0,Gxe0,muxed50);
xor gate_73(Gs1,Gxe1,Gxd1);
xor gate_74(Gs2,muxed66,muxed32);
xor gate_75(Gs3,Gxe3,muxed100);
xor gate_76(Gs4,Gxe4,muxed10);
xor gate_77(Gs5,Gxe5,Gxd5);
xor gate_78(Gs6,muxed14,muxed70);
xor gate_79(Gs7,Gxe7,Gxd7);
not gate_80(Gy0a,Gs0);
not gate_81(Gy1a,Gs1);
not gate_82(Gy2a,muxed42);
not gate_83(Gy0b,Gs0);
not gate_84(Gy1b,Gs1);
not gate_85(Gy3b,Gs3);
not gate_86(Gy0c,Gs0);
not gate_87(Gy2c,muxed42);
not gate_88(Gy3c,Gs3);
not gate_89(Gy1d,Gs1);
not gate_90(Gy2d,muxed42);
not gate_91(Gy3d,Gs3);
not gate_92(Gy5i,Gs5);
not gate_93(Gy7i,Gs7);
not gate_94(Gy5j,Gs5);
not gate_95(Gy6j,muxed91);
not gate_96(Gy4k,muxed49);
not gate_97(Gy7k,Gs7);
not gate_98(Gy4l,muxed49);
not gate_99(Gy6l,muxed91);
not gate_100(Gy4a,muxed49);
not gate_101(Gy5a,Gs5);
not gate_102(Gy6a,muxed91);
not gate_103(Gy4b,muxed49);
not gate_104(Gy5b,Gs5);
not gate_105(Gy7b,Gs7);
not gate_106(Gy4c,muxed49);
not gate_107(Gy6c,muxed91);
not gate_108(Gy7c,Gs7);
not gate_109(Gy5d,Gs5);
not gate_110(Gy6d,muxed91);
not gate_111(Gy7d,Gs7);
not gate_112(Gy1i,Gs1);
not gate_113(Gy3i,Gs3);
not gate_114(Gy1j,Gs1);
not gate_115(Gy2j,muxed42);
not gate_116(Gy0k,Gs0);
not gate_117(Gy3k,Gs3);
not gate_118(Gy0l,Gs0);
not gate_119(Gy2l,muxed42);
and gate_120(Gt0,Gy0a,muxed61,Gy2a,Gs3);
and gate_121(Gt1,Gy0b,Gy1b,muxed42,Gy3b);
and gate_122(Gt2,Gy0c,Gs1,muxed85,Gy3c);
and gate_123(Gt3,Gs0,muxed65,Gy2d,Gy3d);
and gate_124(Gt4,Gy4a,Gy5a,Gy6a,Gs7);
and gate_125(Gt5,Gy4b,Gy5b,muxed91,Gy7b);
and gate_126(Gt6,Gy4c,Gs5,Gy6c,Gy7c);
and gate_127(Gt7,muxed49,Gy5d,muxed102,Gy7d);
or gate_128(Gu0,Gt0,Gt1,Gt2,Gt3);
or gate_129(Gu1,Gt4,muxed71,Gt6,muxed7);
and gate_130(Gwa,muxed49,Gy5i,muxed91,Gy7i,Gu0);
and gate_131(Gwb,muxed49,muxed88,Gy6j,Gs7,Gu0);
and gate_132(Gwc,Gy4k,Gs5,muxed91,Gy7k,Gu0);
and gate_133(Gwd,muxed56,Gs5,muxed99,Gs7,Gu0);
and gate_134(Gwe,Gs0,Gy1i,muxed42,Gy3i,muxed20);
and gate_135(Gwf,Gs0,Gy1j,muxed52,Gs3,muxed20);
and gate_136(Gwg,Gy0k,Gs1,muxed42,Gy3k,muxed20);
and gate_137(Gwh,Gy0l,Gs1,Gy2l,Gs3,muxed20);
and gate_138(Ge0,Gs0,Gwa);
and gate_139(Ge1,Gs1,Gwa);
and gate_140(Ge2,muxed42,Gwa);
and gate_141(Ge3,Gs3,Gwa);
and gate_142(Ge4,Gs0,muxed48);
and gate_143(Ge5,Gs1,muxed48);
and gate_144(Ge6,muxed42,muxed48);
and gate_145(Ge7,Gs3,muxed48);
and gate_146(Ge8,Gs0,Gwc);
and gate_147(Ge9,Gs1,Gwc);
and gate_148(Ge10,muxed42,Gwc);
and gate_149(Ge11,Gs3,Gwc);
and gate_150(Ge12,Gs0,muxed95);
and gate_151(Ge13,Gs1,muxed95);
and gate_152(Ge14,muxed42,muxed95);
and gate_153(Ge15,Gs3,muxed95);
and gate_154(Ge16,muxed49,Gwe);
and gate_155(Ge17,Gs5,Gwe);
and gate_156(Ge18,muxed91,Gwe);
and gate_157(Ge19,Gs7,Gwe);
and gate_158(Ge20,muxed49,muxed73);
and gate_159(Ge21,Gs5,muxed73);
and gate_160(Ge22,muxed91,muxed73);
and gate_161(Ge23,Gs7,muxed73);
and gate_162(Ge24,muxed49,Gwg);
and gate_163(Ge25,Gs5,Gwg);
and gate_164(Ge26,muxed91,Gwg);
and gate_165(Ge27,Gs7,Gwg);
and gate_166(Ge28,muxed49,muxed17);
and gate_167(Ge29,Gs5,muxed17);
and gate_168(Ge30,muxed91,muxed17);
and gate_169(Ge31,Gs7,muxed17);
xor gate_170(God0,Gid0,Ge0);
xor gate_171(God1,Gid1,Ge1);
xor gate_172(God2,Gid2,muxed30);
xor gate_173(God3,Gid3,Ge3);
xor gate_174(God4,Gid4,Ge4);
xor gate_175(God5,Gid5,muxed24);
xor gate_176(God6,Gid6,Ge6);
xor gate_177(God7,Gid7,Ge7);
xor gate_178(God8,Gid8,Ge8);
xor gate_179(God9,Gid9,Ge9);
xor gate_180(God10,Gid10,Ge10);
xor gate_181(God11,Gid11,Ge11);
xor gate_182(God12,Gid12,Ge12);
xor gate_183(God13,Gid13,Ge13);
xor gate_184(God14,Gid14,muxed94);
xor gate_185(God15,Gid15,Ge15);
xor gate_186(God16,Gid16,Ge16);
xor gate_187(God17,Gid17,muxed82);
xor gate_188(God18,Gid18,Ge18);
xor gate_189(God19,Gid19,Ge19);
xor gate_190(God20,Gid20,Ge20);
xor gate_191(God21,Gid21,Ge21);
xor gate_192(God22,Gid22,Ge22);
xor gate_193(God23,Gid23,Ge23);
xor gate_194(God24,muxed53,Ge24);
xor gate_195(God25,Gid25,Ge25);
xor gate_196(God26,Gid26,muxed63);
xor gate_197(God27,Gid27,Ge27);
xor gate_198(God28,Gid28,Ge28);
xor gate_199(God29,Gid29,Ge29);
xor gate_200(God30,Gid30,Ge30);
xor gate_201(God31,Gid31,muxed3);
assign muxed0 = keyinput0 ? Gic4 : muxed1;
assign muxed1 = keyinput1 ? God31 : Gxb1;
assign muxed2 = keyinput2 ? muxed36 : God31;
assign muxed3 = keyinput3 ? muxed16 : Gy7k;
assign muxed4 = keyinput4 ? Gxa5 : muxed16;
assign muxed5 = keyinput5 ? muxed18 : muxed13;
assign muxed6 = keyinput6 ? muxed21 : Gy0k;
assign muxed7 = keyinput7 ? muxed101 : Gh2;
assign muxed8 = keyinput8 ? Gy6l : muxed101;
assign muxed9 = keyinput9 ? Gs4 : muxed50;
assign muxed10 = keyinput10 ? muxed90 : Gy1j;
assign muxed11 = keyinput11 ? Gy5j : muxed90;
assign muxed12 = keyinput12 ? Gh4 : muxed85;
assign muxed13 = keyinput13 ? muxed69 : Gh4;
assign muxed14 = keyinput14 ? Gxe6 : muxed54;
assign muxed15 = keyinput15 ? muxed81 : Gxa15;
assign muxed16 = keyinput16 ? Ge31 : Gt1;
assign muxed17 = keyinput17 ? muxed5 : muxed65;
assign muxed18 = keyinput18 ? Gwh : Ge9;
assign muxed19 = keyinput19 ? muxed46 : Gwh;
assign muxed20 = keyinput20 ? muxed6 : Gy7k;
assign muxed21 = keyinput21 ? muxed89 : muxed92;
assign muxed22 = keyinput22 ? Gy1d : muxed89;
assign muxed23 = keyinput23 ? Gt5 : Gy7i;
assign muxed24 = keyinput24 ? Ge5 : Gt5;
assign muxed25 = keyinput25 ? muxed68 : Gxa11;
assign muxed26 = keyinput26 ? muxed64 : muxed27;
assign muxed27 = keyinput27 ? muxed93 : Ge3;
assign muxed28 = keyinput28 ? Gxa9 : muxed93;
assign muxed29 = keyinput29 ? muxed96 : Ge10;
assign muxed30 = keyinput30 ? Ge2 : muxed96;
assign muxed31 = keyinput31 ? muxed43 : Gs4;
assign muxed32 = keyinput32 ? Gxd2 : Gxc0;
assign muxed33 = keyinput33 ? Gh5 : Gxd2;
assign muxed34 = keyinput34 ? muxed2 : Ge3;
assign muxed35 = keyinput35 ? Gy2j : muxed2;
assign muxed36 = keyinput36 ? muxed45 : Gg7;
assign muxed37 = keyinput37 ? muxed78 : muxed45;
assign muxed38 = keyinput38 ? muxed83 : muxed48;
assign muxed39 = keyinput39 ? Ge17 : muxed83;
assign muxed40 = keyinput40 ? muxed60 : Gy2a;
assign muxed41 = keyinput41 ? Gic0 : muxed42;
assign muxed42 = keyinput42 ? muxed31 : Gs4;
assign muxed43 = keyinput43 ? muxed77 : Gy6l;
assign muxed44 = keyinput44 ? Gxa0 : muxed77;
assign muxed45 = keyinput45 ? muxed19 : Gy7d;
assign muxed46 = keyinput46 ? muxed57 : Gxa2;
assign muxed47 = keyinput47 ? muxed4 : muxed57;
assign muxed48 = keyinput48 ? muxed87 : Gg5;
assign muxed49 = keyinput49 ? muxed9 : Gf5;
assign muxed50 = keyinput50 ? Gxd0 : Gs1;
assign muxed51 = keyinput51 ? Gh0 : muxed20;
assign muxed52 = keyinput52 ? muxed35 : Gh0;
assign muxed53 = keyinput53 ? Gid24 : muxed54;
assign muxed54 = keyinput54 ? muxed15 : Gxa10;
assign muxed55 = keyinput55 ? muxed47 : muxed82;
assign muxed56 = keyinput56 ? Gy4l : muxed47;
assign muxed57 = keyinput57 ? muxed38 : muxed103;
assign muxed58 = keyinput58 ? muxed84 : Gt3;
assign muxed59 = keyinput59 ? muxed40 : muxed87;
assign muxed60 = keyinput60 ? Gf6 : Ge18;
assign muxed61 = keyinput61 ? Gy1a : Gf6;
assign muxed62 = keyinput62 ? muxed26 : Gy3d;
assign muxed63 = keyinput63 ? muxed76 : muxed26;
assign muxed64 = keyinput64 ? Gxa12 : muxed9;
assign muxed65 = keyinput65 ? muxed79 : Gxa12;
assign muxed66 = keyinput66 ? Gxe2 : muxed91;
assign muxed67 = keyinput67 ? muxed25 : Ge30;
assign muxed68 = keyinput68 ? Gs6 : Gy3k;
assign muxed69 = keyinput69 ? Gxa14 : Gs6;
assign muxed70 = keyinput70 ? Gxd6 : Gs3;
assign muxed71 = keyinput71 ? muxed23 : Gxd6;
assign muxed72 = keyinput72 ? Gg2 : Gy2d;
assign muxed73 = keyinput73 ? Gwf : Gg2;
assign muxed74 = keyinput74 ? Gf0 : Gy5b;
assign muxed75 = keyinput75 ? muxed44 : muxed4;
assign muxed76 = keyinput76 ? muxed98 : muxed44;
assign muxed77 = keyinput77 ? muxed37 : Gy3k;
assign muxed78 = keyinput78 ? Gs2 : Gh0;
assign muxed79 = keyinput79 ? muxed22 : Gs2;
assign muxed80 = keyinput80 ? muxed12 : muxed81;
assign muxed81 = keyinput81 ? muxed55 : Gg0;
assign muxed82 = keyinput82 ? muxed39 : Gs5;
assign muxed83 = keyinput83 ? muxed58 : Gg2;
assign muxed84 = keyinput84 ? Gg6 : Gy1i;
assign muxed85 = keyinput85 ? Gy2c : Gg6;
assign muxed86 = keyinput86 ? muxed59 : muxed69;
assign muxed87 = keyinput87 ? Gwb : Gg0;
assign muxed88 = keyinput88 ? muxed11 : Gxd6;
assign muxed89 = keyinput89 ? Gu1 : muxed11;
assign muxed90 = keyinput90 ? Gxd4 : muxed35;
assign muxed91 = keyinput91 ? muxed67 : muxed92;
assign muxed92 = keyinput92 ? muxed28 : muxed79;
assign muxed93 = keyinput93 ? God14 : Gy0l;
assign muxed94 = keyinput94 ? muxed29 : Gxc4;
assign muxed95 = keyinput95 ? muxed97 : muxed29;
assign muxed96 = keyinput96 ? Ge14 : Gy5a;
assign muxed97 = keyinput97 ? Gwd : Gxa6;
assign muxed98 = keyinput98 ? Ge26 : Gwd;
assign muxed99 = keyinput99 ? muxed8 : muxed70;
assign muxed100 = keyinput100 ? Gxd3 : muxed8;
assign muxed101 = keyinput101 ? Gt7 : Gxa10;
assign muxed102 = keyinput102 ? Gy6d : muxed65;
assign muxed103 = keyinput103 ? muxed33 : Gy6d;
endmodule
