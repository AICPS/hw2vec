`timescale 1ns / 1ps
// Verilog
// c432
// Ninputs 36
// Noutputs 7
// NtotalGates 160
// NOT1 40
// NAND2 64
// NOR2 19
// AND9 3
// XOR2 18
// NAND4 14
// AND8 1
// NAND3 1

module top (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
                  N430,N431,N432,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
                  keyinput60, keyinput61, keyinput62, keyinput63,
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
        keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
        keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
        keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
        keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
        keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
                  keyinput134, keyinput135,
        keyinput136, keyinput137, keyinput138, keyinput139, keyinput140,
        keyinput141, keyinput142, keyinput143, keyinput144, keyinput145,
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150,
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155,
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160,
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165,
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170,
        keyinput171);

  input keyinput136, keyinput137, keyinput138, keyinput139, keyinput140;
  input keyinput141, keyinput142, keyinput143, keyinput144, keyinput145;
  input keyinput146, keyinput147, keyinput148, keyinput149, keyinput150;
  input keyinput151, keyinput152, keyinput153, keyinput154, keyinput155;
  input keyinput156, keyinput157, keyinput158, keyinput159, keyinput160;
  input keyinput161, keyinput162, keyinput163, keyinput164, keyinput165;
  input keyinput166, keyinput167, keyinput168, keyinput169, keyinput170;
  input keyinput171;


  input keyinput64, keyinput65, keyinput66, keyinput67, keyinput68;
  input keyinput69, keyinput70, keyinput71, keyinput72, keyinput73;
  input keyinput74, keyinput75, keyinput76, keyinput77, keyinput78;
  input keyinput79, keyinput80, keyinput81, keyinput82, keyinput83;
  input keyinput84, keyinput85, keyinput86, keyinput87, keyinput88;
  input keyinput89, keyinput90, keyinput91, keyinput92, keyinput93;
  input keyinput94, keyinput95, keyinput96, keyinput97, keyinput98;
  input keyinput99, keyinput100, keyinput101, keyinput102, keyinput103;
  input keyinput104, keyinput105, keyinput106, keyinput107, keyinput108;
  input keyinput109, keyinput110, keyinput111, keyinput112, keyinput113;
  input keyinput114, keyinput115, keyinput116, keyinput117, keyinput118;
  input keyinput119, keyinput120, keyinput121, keyinput122, keyinput123;
  input keyinput124, keyinput125, keyinput126, keyinput127, keyinput128;
  input keyinput129, keyinput130, keyinput131, keyinput132, keyinput133;
  input keyinput134, keyinput135;

  wire KeyWire_0_1 , KeyWire_0_2;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31, keyinput32, keyinput33, keyinput34;
  input keyinput35, keyinput36, keyinput37, keyinput38, keyinput39;
  input keyinput40, keyinput41, keyinput42, keyinput43, keyinput44;
  input keyinput45, keyinput46, keyinput47, keyinput48, keyinput49;
  input keyinput50, keyinput51, keyinput52, keyinput53, keyinput54;
  input keyinput55, keyinput56, keyinput57, keyinput58, keyinput59;
  input keyinput60, keyinput61, keyinput62, keyinput63;

  wire [0:63] keyinput_Wire_0;
  wire [0:27] KeyNOTWire_0;

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;

output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429;

not NOT1_1 (N118, N1);
not NOT1_2 (N119, N4);
  not NOT1_3 (keyinput_Wire_0[0], N11);
  xor keyGate_0_0(N122, keyinput0, keyinput_Wire_0[0]);
  not NOT1_4 (keyinput_Wire_0[1], N17);
  xor keyGate_0_1(N123, keyinput1, keyinput_Wire_0[1]);
not NOT1_5 (N126, N24);
not NOT1_6 (N127, N30);
not NOT1_7 (N130, N37);
  not NOT1_8 (keyinput_Wire_0[2], N43);
  xnor keyGate_0_2(N131, keyinput2, keyinput_Wire_0[2]);
  not NOT1_9 (keyinput_Wire_0[3], N50);
  xor keyGate_0_3(N134, keyinput3, keyinput_Wire_0[3]);
not NOT1_10 (N135, N56);
not NOT1_11 (N138, N63);
not NOT1_12 (N139, N69);
  not NOT1_13 (keyinput_Wire_0[4], N76);
  xor keyGate_0_4(KeyNOTWire_0[0], keyinput4, keyinput_Wire_0[4]);
  not KeyNOTGate_0_0(N142, KeyNOTWire_0[0]);
not NOT1_14 (N143, N82);
not NOT1_15 (N146, N89);
not NOT1_16 (N147, N95);
not NOT1_17 (N150, N102);
  not NOT1_18 (keyinput_Wire_0[5], N108);
  xor keyGate_0_5(N151, keyinput5, keyinput_Wire_0[5]);
nand NAND2_19 (N154, N118, N4);
nor NOR2_20 (N157, N8, N119);
  nor NOR2_21 (keyinput_Wire_0[6], N14, N119);
  xnor keyGate_0_6(N158, keyinput6, keyinput_Wire_0[6]);
nand NAND2_22 (N159, N122, N17);
  nand NAND2_23 (keyinput_Wire_0[7], N126, N30);
  xor keyGate_0_7(N162, keyinput7, keyinput_Wire_0[7]);
nand NAND2_24 (N165, N130, N43);
nand NAND2_25 (N168, N134, N56);
  nand NAND2_26 (keyinput_Wire_0[8], N138, N69);
  xor keyGate_0_8(N171, keyinput8, keyinput_Wire_0[8]);
nand NAND2_27 (N174, N142, N82);
  nand NAND2_28 (keyinput_Wire_0[9], N146, N95);
  xnor keyGate_0_9(KeyNOTWire_0[1], keyinput9, keyinput_Wire_0[9]);
  not KeyNOTGate_0_1(N177, KeyNOTWire_0[1]);
nand NAND2_29 (N180, N150, N108);
nor NOR2_30 (N183, N21, N123);
nor NOR2_31 (N184, N27, N123);
nor NOR2_32 (N185, N34, N127);
nor NOR2_33 (N186, N40, N127);
  nor NOR2_34 (keyinput_Wire_0[10], N47, N131);
  xnor keyGate_0_10(KeyNOTWire_0[2], keyinput10, keyinput_Wire_0[10]);
  not KeyNOTGate_0_2(N187, KeyNOTWire_0[2]);
nor NOR2_35 (N188, N53, N131);
nor NOR2_36 (N189, N60, N135);
nor NOR2_37 (N190, N66, N135);
  nor NOR2_38 (keyinput_Wire_0[11], N73, N139);
  xor keyGate_0_11(N191, keyinput11, keyinput_Wire_0[11]);
nor NOR2_39 (N192, N79, N139);
nor NOR2_40 (N193, N86, N143);
nor NOR2_41 (N194, N92, N143);
  nor NOR2_42 (keyinput_Wire_0[12], N99, N147);
  xnor keyGate_0_12(KeyNOTWire_0[3], keyinput12, keyinput_Wire_0[12]);
  not KeyNOTGate_0_3(N195, KeyNOTWire_0[3]);
nor NOR2_43 (N196, N105, N147);
  nor NOR2_44 (keyinput_Wire_0[13], N112, N151);
  xor keyGate_0_13(N197, keyinput13, keyinput_Wire_0[13]);
  nor NOR2_45 (keyinput_Wire_0[14], N115, N151);
  xor keyGate_0_14(N198, keyinput14, keyinput_Wire_0[14]);
and AND9_46 (N199, N154, N159, N162, N165, N168, N171, N174, N177, N180);
not NOT1_47 (N203, N199);
  not NOT1_48 (keyinput_Wire_0[15], N199);
  xor keyGate_0_15(N213, keyinput15, keyinput_Wire_0[15]);
not NOT1_49 (N223, N199);
xor XOR2_50 (N224, N203, N154);
  xor XOR2_51 (keyinput_Wire_0[16], N203, N159);
  xnor keyGate_0_16(KeyNOTWire_0[4], keyinput16, keyinput_Wire_0[16]);
  not KeyNOTGate_0_4(N227, KeyNOTWire_0[4]);
xor XOR2_52 (N230, N203, N162);
xor XOR2_53 (N233, N203, N165);
  xor XOR2_54 (keyinput_Wire_0[17], N203, N168);
  xnor keyGate_0_17(KeyNOTWire_0[5], keyinput17, keyinput_Wire_0[17]);
  not KeyNOTGate_0_5(N236, KeyNOTWire_0[5]);
xor XOR2_55 (N239, N203, N171);
nand NAND2_56 (N242, N1, N213);
  xor XOR2_57 (keyinput_Wire_0[18], N203, N174);
  xnor keyGate_0_18(KeyNOTWire_0[6], keyinput18, keyinput_Wire_0[18]);
  not KeyNOTGate_0_6(N243, KeyNOTWire_0[6]);
  nand NAND2_58 (keyinput_Wire_0[19], N213, N11);
  xor keyGate_0_19(N246, keyinput19, keyinput_Wire_0[19]);
xor XOR2_59 (N247, N203, N177);
  nand NAND2_60 (keyinput_Wire_0[20], N213, N24);
  xor keyGate_0_20(KeyNOTWire_0[7], keyinput20, keyinput_Wire_0[20]);
  not KeyNOTGate_0_7(N250, KeyNOTWire_0[7]);
  xor XOR2_61 (keyinput_Wire_0[21], N203, N180);
  xnor keyGate_0_21(N251, keyinput21, keyinput_Wire_0[21]);
nand NAND2_62 (N254, N213, N37);
  nand NAND2_63 (keyinput_Wire_0[22], N213, N50);
  xnor keyGate_0_22(N255, keyinput22, keyinput_Wire_0[22]);
nand NAND2_64 (N256, N213, N63);
nand NAND2_65 (N257, N213, N76);
  nand NAND2_66 (keyinput_Wire_0[23], N213, N89);
  xor keyGate_0_23(N258, keyinput23, keyinput_Wire_0[23]);
  nand NAND2_67 (keyinput_Wire_0[24], N213, N102);
  xnor keyGate_0_24(N259, keyinput24, keyinput_Wire_0[24]);
  nand NAND2_68 (keyinput_Wire_0[25], N224, N157);
  xnor keyGate_0_25(KeyNOTWire_0[8], keyinput25, keyinput_Wire_0[25]);
  not KeyNOTGate_0_8(N260, KeyNOTWire_0[8]);
  nand NAND2_69 (keyinput_Wire_0[26], N224, N158);
  xnor keyGate_0_26(KeyNOTWire_0[9], keyinput26, keyinput_Wire_0[26]);
  not KeyNOTGate_0_9(N263, KeyNOTWire_0[9]);
  nand NAND2_70 (keyinput_Wire_0[27], N227, N183);
  xor keyGate_0_27(KeyNOTWire_0[10], keyinput27, keyinput_Wire_0[27]);
  not KeyNOTGate_0_10(N264, KeyNOTWire_0[10]);
nand NAND2_71 (N267, N230, N185);
nand NAND2_72 (N270, N233, N187);
nand NAND2_73 (N273, N236, N189);
nand NAND2_74 (N276, N239, N191);
  nand NAND2_75 (keyinput_Wire_0[28], N243, N193);
  xnor keyGate_0_28(N279, keyinput28, keyinput_Wire_0[28]);
  nand NAND2_76 (keyinput_Wire_0[29], N247, N195);
  xor keyGate_0_29(N282, keyinput29, keyinput_Wire_0[29]);
  nand NAND2_77 (keyinput_Wire_0[30], N251, N197);
  xor keyGate_0_30(N285, keyinput30, keyinput_Wire_0[30]);
  nand NAND2_78 (keyinput_Wire_0[31], N227, N184);
  xnor keyGate_0_31(KeyNOTWire_0[11], keyinput31, keyinput_Wire_0[31]);
  not KeyNOTGate_0_11(N288, KeyNOTWire_0[11]);
  nand NAND2_79 (keyinput_Wire_0[32], N230, N186);
  xnor keyGate_0_32(N289, keyinput32, keyinput_Wire_0[32]);
nand NAND2_80 (N290, N233, N188);
  nand NAND2_81 (keyinput_Wire_0[33], N236, N190);
  xor keyGate_0_33(KeyNOTWire_0[12], keyinput33, keyinput_Wire_0[33]);
  not KeyNOTGate_0_12(N291, KeyNOTWire_0[12]);
  nand NAND2_82 (keyinput_Wire_0[34], N239, N192);
  xor keyGate_0_34(N292, keyinput34, keyinput_Wire_0[34]);
nand NAND2_83 (N293, N243, N194);
  nand NAND2_84 (keyinput_Wire_0[35], N247, N196);
  xnor keyGate_0_35(N294, keyinput35, keyinput_Wire_0[35]);
nand NAND2_85 (N295, N251, N198);
  and AND9_86 (keyinput_Wire_0[36], N260, N264, N267, N270, N273, N276, N279, N282, N285);
  xor keyGate_0_36(KeyNOTWire_0[13], keyinput36, keyinput_Wire_0[36]);
  not KeyNOTGate_0_13(N296, KeyNOTWire_0[13]);
  not NOT1_87 (keyinput_Wire_0[37], N263);
  xnor keyGate_0_37(KeyNOTWire_0[14], keyinput37, keyinput_Wire_0[37]);
  not KeyNOTGate_0_14(N300, KeyNOTWire_0[14]);
not NOT1_88 (N301, N288);
not NOT1_89 (N302, N289);
  not NOT1_90 (keyinput_Wire_0[38], N290);
  xor keyGate_0_38(KeyNOTWire_0[15], keyinput38, keyinput_Wire_0[38]);
  not KeyNOTGate_0_15(N303, KeyNOTWire_0[15]);
not NOT1_91 (N304, N291);
not NOT1_92 (N305, N292);
  not NOT1_93 (keyinput_Wire_0[39], N293);
  xnor keyGate_0_39(KeyNOTWire_0[16], keyinput39, keyinput_Wire_0[39]);
  not KeyNOTGate_0_16(N306, KeyNOTWire_0[16]);
  not NOT1_94 (keyinput_Wire_0[40], N294);
  xor keyGate_0_40(KeyNOTWire_0[17], keyinput40, keyinput_Wire_0[40]);
  not KeyNOTGate_0_17(N307, KeyNOTWire_0[17]);
not NOT1_95 (N308, N295);
not NOT1_96 (N309, N296);
not NOT1_97 (N319, N296);
not NOT1_98 (N329, N296);
xor XOR2_99 (N330, N309, N260);
  xor XOR2_100 (keyinput_Wire_0[41], N309, N264);
  xor keyGate_0_41(N331, keyinput41, keyinput_Wire_0[41]);
  xor XOR2_101 (keyinput_Wire_0[42], N309, N267);
  xnor keyGate_0_42(N332, keyinput42, keyinput_Wire_0[42]);
xor XOR2_102 (N333, N309, N270);
nand NAND2_103 (N334, N8, N319);
  xor XOR2_104 (keyinput_Wire_0[43], N309, N273);
  xor keyGate_0_43(N335, keyinput43, keyinput_Wire_0[43]);
  nand NAND2_105 (keyinput_Wire_0[44], N319, N21);
  xor keyGate_0_44(KeyNOTWire_0[18], keyinput44, keyinput_Wire_0[44]);
  not KeyNOTGate_0_18(N336, KeyNOTWire_0[18]);
xor XOR2_106 (N337, N309, N276);
nand NAND2_107 (N338, N319, N34);
xor XOR2_108 (N339, N309, N279);
nand NAND2_109 (N340, N319, N47);
xor XOR2_110 (N341, N309, N282);
nand NAND2_111 (N342, N319, N60);
  xor XOR2_112 (keyinput_Wire_0[45], N309, N285);
  xor keyGate_0_45(KeyNOTWire_0[19], keyinput45, keyinput_Wire_0[45]);
  not KeyNOTGate_0_19(N343, KeyNOTWire_0[19]);
nand NAND2_113 (N344, N319, N73);
nand NAND2_114 (N345, N319, N86);
  nand NAND2_115 (keyinput_Wire_0[46], N319, N99);
  xnor keyGate_0_46(KeyNOTWire_0[20], keyinput46, keyinput_Wire_0[46]);
  not KeyNOTGate_0_20(N346, KeyNOTWire_0[20]);
  nand NAND2_116 (keyinput_Wire_0[47], N319, N112);
  xor keyGate_0_47(N347, keyinput47, keyinput_Wire_0[47]);
nand NAND2_117 (N348, N330, N300);
  nand NAND2_118 (keyinput_Wire_0[48], N331, N301);
  xnor keyGate_0_48(N349, keyinput48, keyinput_Wire_0[48]);
  nand NAND2_119 (keyinput_Wire_0[49], N332, N302);
  xor keyGate_0_49(KeyNOTWire_0[21], keyinput49, keyinput_Wire_0[49]);
  not KeyNOTGate_0_21(N350, KeyNOTWire_0[21]);
nand NAND2_120 (N351, N333, N303);
  nand NAND2_121 (keyinput_Wire_0[50], N335, N304);
  xor keyGate_0_50(N352, keyinput50, keyinput_Wire_0[50]);
  nand NAND2_122 (keyinput_Wire_0[51], N337, N305);
  xnor keyGate_0_51(KeyNOTWire_0[22], keyinput51, keyinput_Wire_0[51]);
  not KeyNOTGate_0_22(N353, KeyNOTWire_0[22]);
  nand NAND2_123 (keyinput_Wire_0[52], N339, N306);
  xnor keyGate_0_52(N354, keyinput52, keyinput_Wire_0[52]);
nand NAND2_124 (N355, N341, N307);
  nand NAND2_125 (keyinput_Wire_0[53], N343, N308);
  xnor keyGate_0_53(N356, keyinput53, keyinput_Wire_0[53]);
and AND9_126 (N357, N348, N349, N350, N351, N352, N353, N354, N355, N356);
not NOT1_127 (N360, N357);
not NOT1_128 (N370, N357);
nand NAND2_129 (N371, N14, N360);
nand NAND2_130 (N372, N360, N27);
  nand NAND2_131 (keyinput_Wire_0[54], N360, N40);
  xnor keyGate_0_54(N373, keyinput54, keyinput_Wire_0[54]);
  nand NAND2_132 (keyinput_Wire_0[55], N360, N53);
  xor keyGate_0_55(KeyNOTWire_0[23], keyinput55, keyinput_Wire_0[55]);
  not KeyNOTGate_0_23(N374, KeyNOTWire_0[23]);
nand NAND2_133 (N375, N360, N66);
  nand NAND2_134 (keyinput_Wire_0[56], N360, N79);
  xnor keyGate_0_56(N376, keyinput56, keyinput_Wire_0[56]);
nand NAND2_135 (N377, N360, N92);
  nand NAND2_136 (keyinput_Wire_0[57], N360, N105);
  xor keyGate_0_57(KeyNOTWire_0[24], keyinput57, keyinput_Wire_0[57]);
  not KeyNOTGate_0_24(N378, KeyNOTWire_0[24]);
  nand NAND2_137 (keyinput_Wire_0[58], N360, N115);
  xnor keyGate_0_58(N379, keyinput58, keyinput_Wire_0[58]);
nand NAND4_138 (N380, N4, N242, N334, N371);
nand NAND4_139 (N381, N246, N336, N372, N17);
  nand NAND4_140 (keyinput_Wire_0[59], N250, N338, N373, N30);
  xor keyGate_0_59(KeyNOTWire_0[25], keyinput59, keyinput_Wire_0[59]);
  not KeyNOTGate_0_25(N386, KeyNOTWire_0[25]);
  nand NAND4_141 (keyinput_Wire_0[60], N254, N340, N374, N43);
  xor keyGate_0_60(N393, keyinput60, keyinput_Wire_0[60]);
nand NAND4_142 (N399, N255, N342, N375, N56);
nand NAND4_143 (N404, N256, N344, N376, N69);
  nand NAND4_144 (keyinput_Wire_0[61], N257, N345, N377, N82);
  xor keyGate_0_61(KeyNOTWire_0[26], keyinput61, keyinput_Wire_0[61]);
  not KeyNOTGate_0_26(N407, KeyNOTWire_0[26]);
nand NAND4_145 (N411, N258, N346, N378, N95);
nand NAND4_146 (N414, N259, N347, N379, N108);
  not NOT1_147 (keyinput_Wire_0[62], N380);
  xnor keyGate_0_62(KeyNOTWire_0[27], keyinput62, keyinput_Wire_0[62]);
  not KeyNOTGate_0_27(N415, KeyNOTWire_0[27]);
and AND8_148 (N416, N381, N386, N393, N399, N404, N407, N411, N414);
not NOT1_149 (N417, N393);
not NOT1_150 (N418, N404);
not NOT1_151 (N419, N407);
not NOT1_152 (N420, N411);
nor NOR2_153 (KeyWire_0_1, N415, N416);
  xor flip_it (N421, KeyWire_0_1, KeyWire_0_2 );
  nand NAND2_154 (keyinput_Wire_0[63], N386, N417);
  xnor keyGate_0_63(N422, keyinput63, keyinput_Wire_0[63]);
nand NAND4_155 (N425, N386, N393, N418, N399);
nand NAND3_156 (N428, N399, N393, N419);
nand NAND4_157 (N429, N386, N393, N407, N420);
nand NAND4_158 (N430, N381, N386, N422, N399);
nand NAND4_159 (N431, N381, N386, N425, N428);
nand NAND4_160 (N432, N381, N422, N425, N429);

AntiSAT some_name( KeyWire_0_2, N17, N86, N4, N21, N8, N76, N47, N102, N53, N108, N82, N79, N73, N50, N92, N11, N105, N63, N37, N27, N56, N66, N115, N99, N69, N24, N112, N14, N30, N95, N89, N40, N34, N1, N60, N43, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135,
       keyinput136, keyinput137, keyinput138, keyinput139, keyinput140,
       keyinput141, keyinput142, keyinput143, keyinput144, keyinput145,
       keyinput146, keyinput147, keyinput148, keyinput149, keyinput150,
       keyinput151, keyinput152, keyinput153, keyinput154, keyinput155,
       keyinput156, keyinput157, keyinput158, keyinput159, keyinput160,
       keyinput161, keyinput162, keyinput163, keyinput164, keyinput165,
       keyinput166, keyinput167, keyinput168, keyinput169, keyinput170,
       keyinput171);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N17, N86, N4, N21, N8, N76, N47, N102, N53, N108, N82, N79, N73, N50, N92, N11, N105, N63, N37, N27, N56, N66, N115, N99, N69, N24, N112, N14, N30, N95, N89, N40, N34, N1, N60, N43, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135 ,
        keyinput136, keyinput137, keyinput138, keyinput139, keyinput140,
        keyinput141, keyinput142, keyinput143, keyinput144, keyinput145,
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150,
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155,
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160,
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165,
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170,
        keyinput171);

  input keyinput136, keyinput137, keyinput138, keyinput139, keyinput140;
  input keyinput141, keyinput142, keyinput143, keyinput144, keyinput145;
  input keyinput146, keyinput147, keyinput148, keyinput149, keyinput150;
  input keyinput151, keyinput152, keyinput153, keyinput154, keyinput155;
  input keyinput156, keyinput157, keyinput158, keyinput159, keyinput160;
  input keyinput161, keyinput162, keyinput163, keyinput164, keyinput165;
  input keyinput166, keyinput167, keyinput168, keyinput169, keyinput170;
  input keyinput171;

  wire [0:35] keyNTin_Wire_1;
  wire [0:15] KeyNOTWire_1;

  input N17, N86, N4, N21, N8, N76, N47, N102, N53, N108, N82, N79, N73, N50, N92, N11, N105, N63, N37, N27, N56, N66, N115, N99, N69, N24, N112, N14, N30, N95, N89, N40, N34, N1, N60, N43;
  input keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73 ;

  xor  KeyGate0 (keyNTin_Wire_1[0], N17, keyinput64);
  xnor keyNTinGate_1_0(newWire_0, keyinput136, keyNTin_Wire_1[0]);
  xnor KeyGate1 (keyNTin_Wire_1[1], N86, keyinput65);
  xnor keyNTinGate_1_1(KeyNOTWire_1[0], keyinput137, keyNTin_Wire_1[1]);
  not KeyNOTGate_1_0(newWire_1, KeyNOTWire_1[0]);
  xnor KeyGate2 (keyNTin_Wire_1[2], N4, keyinput66);
  xor keyNTinGate_1_2(KeyNOTWire_1[1], keyinput138, keyNTin_Wire_1[2]);
  not KeyNOTGate_1_1(newWire_2, KeyNOTWire_1[1]);
  xnor KeyGate3 (newWire_3, N21, keyinput67);
  xor  KeyGate4 (newWire_4, N8, keyinput68);
  xnor KeyGate5 (newWire_5, N76, keyinput69);
  xnor KeyGate6 (newWire_6, N47, keyinput70);
  xnor KeyGate7 (keyNTin_Wire_1[3], N102, keyinput71);
  xnor keyNTinGate_1_3(KeyNOTWire_1[2], keyinput139, keyNTin_Wire_1[3]);
  not KeyNOTGate_1_2(newWire_7, KeyNOTWire_1[2]);
  xor  KeyGate8 (newWire_8, N53, keyinput72);
  xnor KeyGate9 (keyNTin_Wire_1[4], N108, keyinput73);
  xnor keyNTinGate_1_4(newWire_9, keyinput140, keyNTin_Wire_1[4]);
  xor  KeyGate10 (keyNTin_Wire_1[5], N82, keyinput74);
  xor keyNTinGate_1_5(KeyNOTWire_1[3], keyinput141, keyNTin_Wire_1[5]);
  not KeyNOTGate_1_3(newWire_10, KeyNOTWire_1[3]);
  xnor KeyGate11 (keyNTin_Wire_1[6], N79, keyinput75);
  xor keyNTinGate_1_6(newWire_11, keyinput142, keyNTin_Wire_1[6]);
  xor  KeyGate12 (keyNTin_Wire_1[7], N73, keyinput76);
  xnor keyNTinGate_1_7(newWire_12, keyinput143, keyNTin_Wire_1[7]);
  xnor KeyGate13 (newWire_13, N50, keyinput77);
  xnor KeyGate14 (keyNTin_Wire_1[8], N92, keyinput78);
  xnor keyNTinGate_1_8(newWire_14, keyinput144, keyNTin_Wire_1[8]);
  xor  KeyGate15 (newWire_15, N11, keyinput79);
  xor  KeyGate16 (keyNTin_Wire_1[9], N105, keyinput80);
  xnor keyNTinGate_1_9(newWire_16, keyinput145, keyNTin_Wire_1[9]);
  xnor KeyGate17 (newWire_17, N63, keyinput81);
  xnor KeyGate18 (newWire_18, N37, keyinput82);
  xor  KeyGate19 (keyNTin_Wire_1[10], N27, keyinput83);
  xor keyNTinGate_1_10(KeyNOTWire_1[4], keyinput146, keyNTin_Wire_1[10]);
  not KeyNOTGate_1_4(newWire_19, KeyNOTWire_1[4]);
  xor  KeyGate20 (newWire_20, N56, keyinput84);
  xor  KeyGate21 (keyNTin_Wire_1[11], N66, keyinput85);
  xor keyNTinGate_1_11(newWire_21, keyinput147, keyNTin_Wire_1[11]);
  xnor KeyGate22 (keyNTin_Wire_1[12], N115, keyinput86);
  xor keyNTinGate_1_12(newWire_22, keyinput148, keyNTin_Wire_1[12]);
  xnor KeyGate23 (newWire_23, N99, keyinput87);
  xor  KeyGate24 (newWire_24, N69, keyinput88);
  xnor KeyGate25 (newWire_25, N24, keyinput89);
  xnor KeyGate26 (keyNTin_Wire_1[13], N112, keyinput90);
  xnor keyNTinGate_1_13(newWire_26, keyinput149, keyNTin_Wire_1[13]);
  xnor KeyGate27 (newWire_27, N14, keyinput91);
  xnor KeyGate28 (keyNTin_Wire_1[14], N30, keyinput92);
  xor keyNTinGate_1_14(KeyNOTWire_1[5], keyinput150, keyNTin_Wire_1[14]);
  not KeyNOTGate_1_5(newWire_28, KeyNOTWire_1[5]);
  xnor KeyGate29 (keyNTin_Wire_1[15], N95, keyinput93);
  xor keyNTinGate_1_15(KeyNOTWire_1[6], keyinput151, keyNTin_Wire_1[15]);
  not KeyNOTGate_1_6(newWire_29, KeyNOTWire_1[6]);
  xor  KeyGate30 (keyNTin_Wire_1[16], N89, keyinput94);
  xnor keyNTinGate_1_16(newWire_30, keyinput152, keyNTin_Wire_1[16]);
  xnor KeyGate31 (newWire_31, N40, keyinput95);
  xnor KeyGate32 (newWire_32, N34, keyinput96);
  xnor KeyGate33 (keyNTin_Wire_1[17], N1, keyinput97);
  xnor keyNTinGate_1_17(KeyNOTWire_1[7], keyinput153, keyNTin_Wire_1[17]);
  not KeyNOTGate_1_7(newWire_33, KeyNOTWire_1[7]);
  xor  KeyGate34 (newWire_34, N60, keyinput98);
  xor  KeyGate35 (newWire_35, N43, keyinput99);
  xor  KeyGate36 (keyNTin_Wire_1[18], N17, keyinput100);
  xor keyNTinGate_1_18(KeyNOTWire_1[8], keyinput154, keyNTin_Wire_1[18]);
  not KeyNOTGate_1_8(newWire_36, KeyNOTWire_1[8]);
  xor  KeyGate37 (newWire_37, N86, keyinput101);
  xor  KeyGate38 (newWire_38, N4, keyinput102);
  xnor KeyGate39 (newWire_39, N21, keyinput103);
  xnor KeyGate40 (keyNTin_Wire_1[19], N8, keyinput104);
  xnor keyNTinGate_1_19(KeyNOTWire_1[9], keyinput155, keyNTin_Wire_1[19]);
  not KeyNOTGate_1_9(newWire_40, KeyNOTWire_1[9]);
  xor  KeyGate41 (keyNTin_Wire_1[20], N76, keyinput105);
  xnor keyNTinGate_1_20(newWire_41, keyinput156, keyNTin_Wire_1[20]);
  xor  KeyGate42 (keyNTin_Wire_1[21], N47, keyinput106);
  xnor keyNTinGate_1_21(KeyNOTWire_1[10], keyinput157, keyNTin_Wire_1[21]);
  not KeyNOTGate_1_10(newWire_42, KeyNOTWire_1[10]);
  xnor KeyGate43 (newWire_43, N102, keyinput107);
  xor  KeyGate44 (newWire_44, N53, keyinput108);
  xnor KeyGate45 (newWire_45, N108, keyinput109);
  xor  KeyGate46 (keyNTin_Wire_1[22], N82, keyinput110);
  xor keyNTinGate_1_22(newWire_46, keyinput158, keyNTin_Wire_1[22]);
  xnor KeyGate47 (keyNTin_Wire_1[23], N79, keyinput111);
  xnor keyNTinGate_1_23(KeyNOTWire_1[11], keyinput159, keyNTin_Wire_1[23]);
  not KeyNOTGate_1_11(newWire_47, KeyNOTWire_1[11]);
  xnor KeyGate48 (keyNTin_Wire_1[24], N73, keyinput112);
  xor keyNTinGate_1_24(newWire_48, keyinput160, keyNTin_Wire_1[24]);
  xor  KeyGate49 (newWire_49, N50, keyinput113);
  xnor KeyGate50 (newWire_50, N92, keyinput114);
  xnor KeyGate51 (newWire_51, N11, keyinput115);
  xor  KeyGate52 (keyNTin_Wire_1[25], N105, keyinput116);
  xnor keyNTinGate_1_25(KeyNOTWire_1[12], keyinput161, keyNTin_Wire_1[25]);
  not KeyNOTGate_1_12(newWire_52, KeyNOTWire_1[12]);
  xnor KeyGate53 (newWire_53, N63, keyinput117);
  xor  KeyGate54 (keyNTin_Wire_1[26], N37, keyinput118);
  xor keyNTinGate_1_26(newWire_54, keyinput162, keyNTin_Wire_1[26]);
  xnor KeyGate55 (newWire_55, N27, keyinput119);
  xor  KeyGate56 (newWire_56, N56, keyinput120);
  xnor KeyGate57 (newWire_57, N66, keyinput121);
  xnor KeyGate58 (keyNTin_Wire_1[27], N115, keyinput122);
  xnor keyNTinGate_1_27(newWire_58, keyinput163, keyNTin_Wire_1[27]);
  xor  KeyGate59 (keyNTin_Wire_1[28], N99, keyinput123);
  xor keyNTinGate_1_28(newWire_59, keyinput164, keyNTin_Wire_1[28]);
  xor  KeyGate60 (keyNTin_Wire_1[29], N69, keyinput124);
  xor keyNTinGate_1_29(newWire_60, keyinput165, keyNTin_Wire_1[29]);
  xnor KeyGate61 (keyNTin_Wire_1[30], N24, keyinput125);
  xnor keyNTinGate_1_30(KeyNOTWire_1[13], keyinput166, keyNTin_Wire_1[30]);
  not KeyNOTGate_1_13(newWire_61, KeyNOTWire_1[13]);
  xnor KeyGate62 (keyNTin_Wire_1[31], N112, keyinput126);
  xor keyNTinGate_1_31(newWire_62, keyinput167, keyNTin_Wire_1[31]);
  xor  KeyGate63 (newWire_63, N14, keyinput127);
  xnor KeyGate64 (keyNTin_Wire_1[32], N30, keyinput128);
  xnor keyNTinGate_1_32(newWire_64, keyinput168, keyNTin_Wire_1[32]);
  xnor KeyGate65 (newWire_65, N95, keyinput129);
  xor  KeyGate66 (newWire_66, N89, keyinput130);
  xor  KeyGate67 (keyNTin_Wire_1[33], N40, keyinput131);
  xnor keyNTinGate_1_33(KeyNOTWire_1[14], keyinput169, keyNTin_Wire_1[33]);
  not KeyNOTGate_1_14(newWire_67, KeyNOTWire_1[14]);
  xnor KeyGate68 (keyNTin_Wire_1[34], N34, keyinput132);
  xnor keyNTinGate_1_34(newWire_68, keyinput170, keyNTin_Wire_1[34]);
  xor  KeyGate69 (newWire_69, N1, keyinput133);
  xnor KeyGate70 (keyNTin_Wire_1[35], N60, keyinput134);
  xor keyNTinGate_1_35(KeyNOTWire_1[15], keyinput171, keyNTin_Wire_1[35]);
  not KeyNOTGate_1_15(newWire_70, KeyNOTWire_1[15]);
  xnor KeyGate71 (newWire_71, N43, keyinput135);
  and some_function (newWire_72, newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35 );
  nand compl_function (newWire_73, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71);
  and finalAND (KeyWire_0_2, newWire_72, newWire_73);

endmodule /* AntiSAT */
