`timescale 1ns / 1ps
// Verilog
// c880
// Ninputs 60
// Noutputs 26
// NtotalGates 383
// NAND4 13
// AND3 12
// NAND2 60
// NAND3 14
// AND2 105
// OR2 29
// NOT1 63
// NOR2 61
// BUFF1 26

module top (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
                  N865,N866,N874,N878,N879,N880,
        keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4,
        keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9,
        keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14,
        keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19,
        keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24,
        keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29,
        keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34,
        keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39,
        keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44,
        keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49,
        keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54,
        keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59,
        keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64,
        keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69,
        keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74,
        keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79,
        keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84,
        keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89,
        keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94,
        keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99,
        keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104,
        keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109,
        keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114,
        keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119,
        keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124,
        keyIn_0_125, keyIn_0_126, keyIn_0_127);

  input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4;
  input keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9;
  input keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14;
  input keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19;
  input keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24;
  input keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29;
  input keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34;
  input keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39;
  input keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44;
  input keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49;
  input keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54;
  input keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59;
  input keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64;
  input keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69;
  input keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74;
  input keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79;
  input keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84;
  input keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89;
  input keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94;
  input keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99;
  input keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104;
  input keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109;
  input keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114;
  input keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119;
  input keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124;
  input keyIn_0_125, keyIn_0_126, keyIn_0_127;

  wire [0:127] KeyWire_0;
  wire [0:63] KeyNOTWire_0;

input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;

output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;

wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877;

nand NAND4_1 (N269, N1, N8, N13, N17);
nand NAND4_2 (N270, N1, N26, N13, N17);
and AND3_3 (N273, N29, N36, N42);
  and AND3_4 (KeyWire_0[0], N1, N26, N51);
  xnor KeyGate_0_0(KeyNOTWire_0[0], keyIn_0_0, KeyWire_0[0]);
  not KeyNOTGate_0_0(N276, KeyNOTWire_0[0]);
  nand NAND4_5 (KeyWire_0[1], N1, N8, N51, N17);
  xnor KeyGate_0_1(N279, keyIn_0_1, KeyWire_0[1]);
nand NAND4_6 (N280, N1, N8, N13, N55);
nand NAND4_7 (N284, N59, N42, N68, N72);
nand NAND2_8 (N285, N29, N68);
nand NAND3_9 (N286, N59, N68, N74);
  and AND3_10 (KeyWire_0[2], N29, N75, N80);
  xor KeyGate_0_2(KeyNOTWire_0[1], keyIn_0_2, KeyWire_0[2]);
  not KeyNOTGate_0_1(N287, KeyNOTWire_0[1]);
and AND3_11 (N290, N29, N75, N42);
and AND3_12 (N291, N29, N36, N80);
and AND3_13 (N292, N29, N36, N42);
and AND3_14 (N293, N59, N75, N80);
  and AND3_15 (KeyWire_0[3], N59, N75, N42);
  xnor KeyGate_0_3(KeyNOTWire_0[2], keyIn_0_3, KeyWire_0[3]);
  not KeyNOTGate_0_2(N294, KeyNOTWire_0[2]);
and AND3_16 (N295, N59, N36, N80);
and AND3_17 (N296, N59, N36, N42);
and AND2_18 (N297, N85, N86);
or OR2_19 (N298, N87, N88);
nand NAND2_20 (N301, N91, N96);
or OR2_21 (N302, N91, N96);
nand NAND2_22 (N303, N101, N106);
or OR2_23 (N304, N101, N106);
nand NAND2_24 (N305, N111, N116);
or OR2_25 (N306, N111, N116);
nand NAND2_26 (N307, N121, N126);
or OR2_27 (N308, N121, N126);
and AND2_28 (N309, N8, N138);
  not NOT1_29 (KeyWire_0[4], N268);
  xor KeyGate_0_4(KeyNOTWire_0[3], keyIn_0_4, KeyWire_0[4]);
  not KeyNOTGate_0_3(N310, KeyNOTWire_0[3]);
and AND2_30 (N316, N51, N138);
and AND2_31 (N317, N17, N138);
and AND2_32 (N318, N152, N138);
  nand NAND2_33 (KeyWire_0[5], N59, N156);
  xor KeyGate_0_5(KeyNOTWire_0[4], keyIn_0_5, KeyWire_0[5]);
  not KeyNOTGate_0_4(N319, KeyNOTWire_0[4]);
  nor NOR2_34 (KeyWire_0[6], N17, N42);
  xor KeyGate_0_6(KeyNOTWire_0[5], keyIn_0_6, KeyWire_0[6]);
  not KeyNOTGate_0_5(N322, KeyNOTWire_0[5]);
  and AND2_35 (KeyWire_0[7], N17, N42);
  xor KeyGate_0_7(N323, keyIn_0_7, KeyWire_0[7]);
nand NAND2_36 (N324, N159, N165);
or OR2_37 (N325, N159, N165);
nand NAND2_38 (N326, N171, N177);
or OR2_39 (N327, N171, N177);
nand NAND2_40 (N328, N183, N189);
or OR2_41 (N329, N183, N189);
nand NAND2_42 (N330, N195, N201);
or OR2_43 (N331, N195, N201);
and AND2_44 (N332, N210, N91);
and AND2_45 (N333, N210, N96);
and AND2_46 (N334, N210, N101);
and AND2_47 (N335, N210, N106);
and AND2_48 (N336, N210, N111);
and AND2_49 (N337, N255, N259);
and AND2_50 (N338, N210, N116);
and AND2_51 (N339, N255, N260);
and AND2_52 (N340, N210, N121);
and AND2_53 (N341, N255, N267);
not NOT1_54 (N342, N269);
not NOT1_55 (N343, N273);
or OR2_56 (N344, N270, N273);
  not NOT1_57 (KeyWire_0[8], N276);
  xnor KeyGate_0_8(N345, keyIn_0_8, KeyWire_0[8]);
not NOT1_58 (N346, N276);
  not NOT1_59 (KeyWire_0[9], N279);
  xor KeyGate_0_9(N347, keyIn_0_9, KeyWire_0[9]);
  nor NOR2_60 (KeyWire_0[10], N280, N284);
  xor KeyGate_0_10(KeyNOTWire_0[6], keyIn_0_10, KeyWire_0[10]);
  not KeyNOTGate_0_6(N348, KeyNOTWire_0[6]);
or OR2_61 (N349, N280, N285);
or OR2_62 (N350, N280, N286);
not NOT1_63 (N351, N293);
  not NOT1_64 (KeyWire_0[11], N294);
  xnor KeyGate_0_11(KeyNOTWire_0[7], keyIn_0_11, KeyWire_0[11]);
  not KeyNOTGate_0_7(N352, KeyNOTWire_0[7]);
not NOT1_65 (N353, N295);
not NOT1_66 (N354, N296);
nand NAND2_67 (N355, N89, N298);
and AND2_68 (N356, N90, N298);
  nand NAND2_69 (KeyWire_0[12], N301, N302);
  xor KeyGate_0_12(N357, keyIn_0_12, KeyWire_0[12]);
  nand NAND2_70 (KeyWire_0[13], N303, N304);
  xnor KeyGate_0_13(KeyNOTWire_0[8], keyIn_0_13, KeyWire_0[13]);
  not KeyNOTGate_0_8(N360, KeyNOTWire_0[8]);
  nand NAND2_71 (KeyWire_0[14], N305, N306);
  xnor KeyGate_0_14(KeyNOTWire_0[9], keyIn_0_14, KeyWire_0[14]);
  not KeyNOTGate_0_9(N363, KeyNOTWire_0[9]);
  nand NAND2_72 (KeyWire_0[15], N307, N308);
  xor KeyGate_0_15(N366, keyIn_0_15, KeyWire_0[15]);
  not NOT1_73 (KeyWire_0[16], N310);
  xnor KeyGate_0_16(N369, keyIn_0_16, KeyWire_0[16]);
  nor NOR2_74 (KeyWire_0[17], N322, N323);
  xor KeyGate_0_17(N375, keyIn_0_17, KeyWire_0[17]);
  nand NAND2_75 (KeyWire_0[18], N324, N325);
  xnor KeyGate_0_18(N376, keyIn_0_18, KeyWire_0[18]);
  nand NAND2_76 (KeyWire_0[19], N326, N327);
  xor KeyGate_0_19(N379, keyIn_0_19, KeyWire_0[19]);
  nand NAND2_77 (KeyWire_0[20], N328, N329);
  xor KeyGate_0_20(KeyNOTWire_0[10], keyIn_0_20, KeyWire_0[20]);
  not KeyNOTGate_0_10(N382, KeyNOTWire_0[10]);
  nand NAND2_78 (KeyWire_0[21], N330, N331);
  xnor KeyGate_0_21(KeyNOTWire_0[11], keyIn_0_21, KeyWire_0[21]);
  not KeyNOTGate_0_11(N385, KeyNOTWire_0[11]);
buf BUFF1_79 (N388, N290);
buf BUFF1_80 (N389, N291);
buf BUFF1_81 (N390, N292);
buf BUFF1_82 (N391, N297);
or OR2_83 (N392, N270, N343);
  not NOT1_84 (KeyWire_0[22], N345);
  xor KeyGate_0_22(KeyNOTWire_0[12], keyIn_0_22, KeyWire_0[22]);
  not KeyNOTGate_0_12(N393, KeyNOTWire_0[12]);
not NOT1_85 (N399, N346);
and AND2_86 (N400, N348, N73);
not NOT1_87 (N401, N349);
not NOT1_88 (N402, N350);
not NOT1_89 (N403, N355);
not NOT1_90 (N404, N357);
not NOT1_91 (N405, N360);
  and AND2_92 (KeyWire_0[23], N357, N360);
  xor KeyGate_0_23(N406, keyIn_0_23, KeyWire_0[23]);
not NOT1_93 (N407, N363);
not NOT1_94 (N408, N366);
  and AND2_95 (KeyWire_0[24], N363, N366);
  xor KeyGate_0_24(KeyNOTWire_0[13], keyIn_0_24, KeyWire_0[24]);
  not KeyNOTGate_0_13(N409, KeyNOTWire_0[13]);
  nand NAND2_96 (KeyWire_0[25], N347, N352);
  xnor KeyGate_0_25(KeyNOTWire_0[14], keyIn_0_25, KeyWire_0[25]);
  not KeyNOTGate_0_14(N410, KeyNOTWire_0[14]);
not NOT1_97 (N411, N376);
not NOT1_98 (N412, N379);
  and AND2_99 (KeyWire_0[26], N376, N379);
  xnor KeyGate_0_26(KeyNOTWire_0[15], keyIn_0_26, KeyWire_0[26]);
  not KeyNOTGate_0_15(N413, KeyNOTWire_0[15]);
not NOT1_100 (N414, N382);
not NOT1_101 (N415, N385);
  and AND2_102 (KeyWire_0[27], N382, N385);
  xnor KeyGate_0_27(N416, keyIn_0_27, KeyWire_0[27]);
and AND2_103 (N417, N210, N369);
buf BUFF1_104 (N418, N342);
buf BUFF1_105 (N419, N344);
buf BUFF1_106 (N420, N351);
buf BUFF1_107 (N421, N353);
buf BUFF1_108 (N422, N354);
buf BUFF1_109 (N423, N356);
not NOT1_110 (N424, N400);
  and AND2_111 (KeyWire_0[28], N404, N405);
  xor KeyGate_0_28(N425, keyIn_0_28, KeyWire_0[28]);
  and AND2_112 (KeyWire_0[29], N407, N408);
  xnor KeyGate_0_29(N426, keyIn_0_29, KeyWire_0[29]);
  and AND3_113 (KeyWire_0[30], N319, N393, N55);
  xnor KeyGate_0_30(N427, keyIn_0_30, KeyWire_0[30]);
  and AND3_114 (KeyWire_0[31], N393, N17, N287);
  xnor KeyGate_0_31(N432, keyIn_0_31, KeyWire_0[31]);
  nand NAND3_115 (KeyWire_0[32], N393, N287, N55);
  xnor KeyGate_0_32(KeyNOTWire_0[16], keyIn_0_32, KeyWire_0[32]);
  not KeyNOTGate_0_16(N437, KeyNOTWire_0[16]);
  nand NAND4_116 (KeyWire_0[33], N375, N59, N156, N393);
  xor KeyGate_0_33(KeyNOTWire_0[17], keyIn_0_33, KeyWire_0[33]);
  not KeyNOTGate_0_17(N442, KeyNOTWire_0[17]);
  nand NAND3_117 (KeyWire_0[34], N393, N319, N17);
  xnor KeyGate_0_34(N443, keyIn_0_34, KeyWire_0[34]);
  and AND2_118 (KeyWire_0[35], N411, N412);
  xor KeyGate_0_35(N444, keyIn_0_35, KeyWire_0[35]);
  and AND2_119 (KeyWire_0[36], N414, N415);
  xor KeyGate_0_36(N445, keyIn_0_36, KeyWire_0[36]);
buf BUFF1_120 (N446, N392);
buf BUFF1_121 (N447, N399);
buf BUFF1_122 (N448, N401);
buf BUFF1_123 (N449, N402);
buf BUFF1_124 (N450, N403);
not NOT1_125 (N451, N424);
  nor NOR2_126 (KeyWire_0[37], N406, N425);
  xor KeyGate_0_37(KeyNOTWire_0[18], keyIn_0_37, KeyWire_0[37]);
  not KeyNOTGate_0_18(N460, KeyNOTWire_0[18]);
  nor NOR2_127 (KeyWire_0[38], N409, N426);
  xor KeyGate_0_38(N463, keyIn_0_38, KeyWire_0[38]);
  nand NAND2_128 (KeyWire_0[39], N442, N410);
  xnor KeyGate_0_39(N466, keyIn_0_39, KeyWire_0[39]);
and AND2_129 (N475, N143, N427);
  and AND2_130 (KeyWire_0[40], N310, N432);
  xnor KeyGate_0_40(KeyNOTWire_0[19], keyIn_0_40, KeyWire_0[40]);
  not KeyNOTGate_0_19(N476, KeyNOTWire_0[19]);
and AND2_131 (N477, N146, N427);
  and AND2_132 (KeyWire_0[41], N310, N432);
  xnor KeyGate_0_41(KeyNOTWire_0[20], keyIn_0_41, KeyWire_0[41]);
  not KeyNOTGate_0_20(N478, KeyNOTWire_0[20]);
and AND2_133 (N479, N149, N427);
  and AND2_134 (KeyWire_0[42], N310, N432);
  xor KeyGate_0_42(KeyNOTWire_0[21], keyIn_0_42, KeyWire_0[42]);
  not KeyNOTGate_0_21(N480, KeyNOTWire_0[21]);
and AND2_135 (N481, N153, N427);
  and AND2_136 (KeyWire_0[43], N310, N432);
  xor KeyGate_0_43(KeyNOTWire_0[22], keyIn_0_43, KeyWire_0[43]);
  not KeyNOTGate_0_22(N482, KeyNOTWire_0[22]);
  nand NAND2_137 (KeyWire_0[44], N443, N1);
  xor KeyGate_0_44(N483, keyIn_0_44, KeyWire_0[44]);
  or OR2_138 (KeyWire_0[45], N369, N437);
  xor KeyGate_0_45(KeyNOTWire_0[23], keyIn_0_45, KeyWire_0[45]);
  not KeyNOTGate_0_23(N488, KeyNOTWire_0[23]);
  or OR2_139 (KeyWire_0[46], N369, N437);
  xor KeyGate_0_46(N489, keyIn_0_46, KeyWire_0[46]);
  or OR2_140 (KeyWire_0[47], N369, N437);
  xor KeyGate_0_47(N490, keyIn_0_47, KeyWire_0[47]);
  or OR2_141 (KeyWire_0[48], N369, N437);
  xor KeyGate_0_48(KeyNOTWire_0[24], keyIn_0_48, KeyWire_0[48]);
  not KeyNOTGate_0_24(N491, KeyNOTWire_0[24]);
  nor NOR2_142 (KeyWire_0[49], N413, N444);
  xor KeyGate_0_49(N492, keyIn_0_49, KeyWire_0[49]);
  nor NOR2_143 (KeyWire_0[50], N416, N445);
  xnor KeyGate_0_50(KeyNOTWire_0[25], keyIn_0_50, KeyWire_0[50]);
  not KeyNOTGate_0_25(N495, KeyNOTWire_0[25]);
nand NAND2_144 (N498, N130, N460);
or OR2_145 (N499, N130, N460);
nand NAND2_146 (N500, N463, N135);
or OR2_147 (N501, N463, N135);
and AND2_148 (N502, N91, N466);
  nor NOR2_149 (KeyWire_0[51], N475, N476);
  xnor KeyGate_0_51(KeyNOTWire_0[26], keyIn_0_51, KeyWire_0[51]);
  not KeyNOTGate_0_26(N503, KeyNOTWire_0[26]);
and AND2_150 (N504, N96, N466);
  nor NOR2_151 (KeyWire_0[52], N477, N478);
  xnor KeyGate_0_52(KeyNOTWire_0[27], keyIn_0_52, KeyWire_0[52]);
  not KeyNOTGate_0_27(N505, KeyNOTWire_0[27]);
and AND2_152 (N506, N101, N466);
  nor NOR2_153 (KeyWire_0[53], N479, N480);
  xor KeyGate_0_53(KeyNOTWire_0[28], keyIn_0_53, KeyWire_0[53]);
  not KeyNOTGate_0_28(N507, KeyNOTWire_0[28]);
and AND2_154 (N508, N106, N466);
  nor NOR2_155 (KeyWire_0[54], N481, N482);
  xnor KeyGate_0_54(N509, keyIn_0_54, KeyWire_0[54]);
  and AND2_156 (KeyWire_0[55], N143, N483);
  xor KeyGate_0_55(N510, keyIn_0_55, KeyWire_0[55]);
  and AND2_157 (KeyWire_0[56], N111, N466);
  xor KeyGate_0_56(KeyNOTWire_0[29], keyIn_0_56, KeyWire_0[56]);
  not KeyNOTGate_0_29(N511, KeyNOTWire_0[29]);
  and AND2_158 (KeyWire_0[57], N146, N483);
  xor KeyGate_0_57(N512, keyIn_0_57, KeyWire_0[57]);
  and AND2_159 (KeyWire_0[58], N116, N466);
  xor KeyGate_0_58(KeyNOTWire_0[30], keyIn_0_58, KeyWire_0[58]);
  not KeyNOTGate_0_30(N513, KeyNOTWire_0[30]);
  and AND2_160 (KeyWire_0[59], N149, N483);
  xor KeyGate_0_59(KeyNOTWire_0[31], keyIn_0_59, KeyWire_0[59]);
  not KeyNOTGate_0_31(N514, KeyNOTWire_0[31]);
  and AND2_161 (KeyWire_0[60], N121, N466);
  xor KeyGate_0_60(KeyNOTWire_0[32], keyIn_0_60, KeyWire_0[60]);
  not KeyNOTGate_0_32(N515, KeyNOTWire_0[32]);
  and AND2_162 (KeyWire_0[61], N153, N483);
  xor KeyGate_0_61(N516, keyIn_0_61, KeyWire_0[61]);
  and AND2_163 (KeyWire_0[62], N126, N466);
  xnor KeyGate_0_62(KeyNOTWire_0[33], keyIn_0_62, KeyWire_0[62]);
  not KeyNOTGate_0_33(N517, KeyNOTWire_0[33]);
nand NAND2_164 (N518, N130, N492);
or OR2_165 (N519, N130, N492);
nand NAND2_166 (N520, N495, N207);
or OR2_167 (N521, N495, N207);
and AND2_168 (N522, N451, N159);
and AND2_169 (N523, N451, N165);
and AND2_170 (N524, N451, N171);
and AND2_171 (N525, N451, N177);
and AND2_172 (N526, N451, N183);
nand NAND2_173 (N527, N451, N189);
nand NAND2_174 (N528, N451, N195);
nand NAND2_175 (N529, N451, N201);
nand NAND2_176 (N530, N498, N499);
nand NAND2_177 (N533, N500, N501);
  nor NOR2_178 (KeyWire_0[63], N309, N502);
  xor KeyGate_0_63(KeyNOTWire_0[34], keyIn_0_63, KeyWire_0[63]);
  not KeyNOTGate_0_34(N536, KeyNOTWire_0[34]);
  nor NOR2_179 (KeyWire_0[64], N316, N504);
  xnor KeyGate_0_64(N537, keyIn_0_64, KeyWire_0[64]);
  nor NOR2_180 (KeyWire_0[65], N317, N506);
  xnor KeyGate_0_65(KeyNOTWire_0[35], keyIn_0_65, KeyWire_0[65]);
  not KeyNOTGate_0_35(N538, KeyNOTWire_0[35]);
  nor NOR2_181 (KeyWire_0[66], N318, N508);
  xor KeyGate_0_66(N539, keyIn_0_66, KeyWire_0[66]);
  nor NOR2_182 (KeyWire_0[67], N510, N511);
  xnor KeyGate_0_67(KeyNOTWire_0[36], keyIn_0_67, KeyWire_0[67]);
  not KeyNOTGate_0_36(N540, KeyNOTWire_0[36]);
  nor NOR2_183 (KeyWire_0[68], N512, N513);
  xnor KeyGate_0_68(KeyNOTWire_0[37], keyIn_0_68, KeyWire_0[68]);
  not KeyNOTGate_0_37(N541, KeyNOTWire_0[37]);
  nor NOR2_184 (KeyWire_0[69], N514, N515);
  xnor KeyGate_0_69(N542, keyIn_0_69, KeyWire_0[69]);
  nor NOR2_185 (KeyWire_0[70], N516, N517);
  xor KeyGate_0_70(N543, keyIn_0_70, KeyWire_0[70]);
nand NAND2_186 (N544, N518, N519);
nand NAND2_187 (N547, N520, N521);
not NOT1_188 (N550, N530);
not NOT1_189 (N551, N533);
and AND2_190 (N552, N530, N533);
  nand NAND2_191 (KeyWire_0[71], N536, N503);
  xnor KeyGate_0_71(N553, keyIn_0_71, KeyWire_0[71]);
  nand NAND2_192 (KeyWire_0[72], N537, N505);
  xor KeyGate_0_72(N557, keyIn_0_72, KeyWire_0[72]);
  nand NAND2_193 (KeyWire_0[73], N538, N507);
  xnor KeyGate_0_73(KeyNOTWire_0[38], keyIn_0_73, KeyWire_0[73]);
  not KeyNOTGate_0_38(N561, KeyNOTWire_0[38]);
  nand NAND2_194 (KeyWire_0[74], N539, N509);
  xor KeyGate_0_74(N565, keyIn_0_74, KeyWire_0[74]);
  nand NAND2_195 (KeyWire_0[75], N488, N540);
  xor KeyGate_0_75(N569, keyIn_0_75, KeyWire_0[75]);
  nand NAND2_196 (KeyWire_0[76], N489, N541);
  xor KeyGate_0_76(KeyNOTWire_0[39], keyIn_0_76, KeyWire_0[76]);
  not KeyNOTGate_0_39(N573, KeyNOTWire_0[39]);
  nand NAND2_197 (KeyWire_0[77], N490, N542);
  xnor KeyGate_0_77(N577, keyIn_0_77, KeyWire_0[77]);
  nand NAND2_198 (KeyWire_0[78], N491, N543);
  xnor KeyGate_0_78(N581, keyIn_0_78, KeyWire_0[78]);
not NOT1_199 (N585, N544);
not NOT1_200 (N586, N547);
and AND2_201 (N587, N544, N547);
and AND2_202 (N588, N550, N551);
and AND2_203 (N589, N585, N586);
nand NAND2_204 (N590, N553, N159);
or OR2_205 (N593, N553, N159);
and AND2_206 (N596, N246, N553);
nand NAND2_207 (N597, N557, N165);
or OR2_208 (N600, N557, N165);
and AND2_209 (N605, N246, N557);
nand NAND2_210 (N606, N561, N171);
or OR2_211 (N609, N561, N171);
and AND2_212 (N615, N246, N561);
nand NAND2_213 (N616, N565, N177);
or OR2_214 (N619, N565, N177);
and AND2_215 (N624, N246, N565);
nand NAND2_216 (N625, N569, N183);
or OR2_217 (N628, N569, N183);
and AND2_218 (N631, N246, N569);
  nand NAND2_219 (KeyWire_0[79], N573, N189);
  xor KeyGate_0_79(N632, keyIn_0_79, KeyWire_0[79]);
  or OR2_220 (KeyWire_0[80], N573, N189);
  xor KeyGate_0_80(N635, keyIn_0_80, KeyWire_0[80]);
and AND2_221 (N640, N246, N573);
  nand NAND2_222 (KeyWire_0[81], N577, N195);
  xor KeyGate_0_81(KeyNOTWire_0[40], keyIn_0_81, KeyWire_0[81]);
  not KeyNOTGate_0_40(N641, KeyNOTWire_0[40]);
  or OR2_223 (KeyWire_0[82], N577, N195);
  xnor KeyGate_0_82(N644, keyIn_0_82, KeyWire_0[82]);
and AND2_224 (N650, N246, N577);
  nand NAND2_225 (KeyWire_0[83], N581, N201);
  xnor KeyGate_0_83(N651, keyIn_0_83, KeyWire_0[83]);
  or OR2_226 (KeyWire_0[84], N581, N201);
  xor KeyGate_0_84(KeyNOTWire_0[41], keyIn_0_84, KeyWire_0[84]);
  not KeyNOTGate_0_41(N654, KeyNOTWire_0[41]);
and AND2_227 (N659, N246, N581);
nor NOR2_228 (N660, N552, N588);
nor NOR2_229 (N661, N587, N589);
not NOT1_230 (N662, N590);
  and AND2_231 (KeyWire_0[85], N593, N590);
  xor KeyGate_0_85(KeyNOTWire_0[42], keyIn_0_85, KeyWire_0[85]);
  not KeyNOTGate_0_42(N665, KeyNOTWire_0[42]);
nor NOR2_232 (N669, N596, N522);
not NOT1_233 (N670, N597);
  and AND2_234 (KeyWire_0[86], N600, N597);
  xor KeyGate_0_86(KeyNOTWire_0[43], keyIn_0_86, KeyWire_0[86]);
  not KeyNOTGate_0_43(N673, KeyNOTWire_0[43]);
nor NOR2_235 (N677, N605, N523);
not NOT1_236 (N678, N606);
  and AND2_237 (KeyWire_0[87], N609, N606);
  xnor KeyGate_0_87(N682, keyIn_0_87, KeyWire_0[87]);
nor NOR2_238 (N686, N615, N524);
not NOT1_239 (N687, N616);
  and AND2_240 (KeyWire_0[88], N619, N616);
  xnor KeyGate_0_88(KeyNOTWire_0[44], keyIn_0_88, KeyWire_0[88]);
  not KeyNOTGate_0_44(N692, KeyNOTWire_0[44]);
nor NOR2_241 (N696, N624, N525);
not NOT1_242 (N697, N625);
  and AND2_243 (KeyWire_0[89], N628, N625);
  xnor KeyGate_0_89(N700, keyIn_0_89, KeyWire_0[89]);
nor NOR2_244 (N704, N631, N526);
not NOT1_245 (N705, N632);
  and AND2_246 (KeyWire_0[90], N635, N632);
  xnor KeyGate_0_90(KeyNOTWire_0[45], keyIn_0_90, KeyWire_0[90]);
  not KeyNOTGate_0_45(N708, KeyNOTWire_0[45]);
nor NOR2_247 (N712, N337, N640);
  not NOT1_248 (KeyWire_0[91], N641);
  xor KeyGate_0_91(KeyNOTWire_0[46], keyIn_0_91, KeyWire_0[91]);
  not KeyNOTGate_0_46(N713, KeyNOTWire_0[46]);
  and AND2_249 (KeyWire_0[92], N644, N641);
  xnor KeyGate_0_92(N717, keyIn_0_92, KeyWire_0[92]);
nor NOR2_250 (N721, N339, N650);
  not NOT1_251 (KeyWire_0[93], N651);
  xor KeyGate_0_93(KeyNOTWire_0[47], keyIn_0_93, KeyWire_0[93]);
  not KeyNOTGate_0_47(N722, KeyNOTWire_0[47]);
  and AND2_252 (KeyWire_0[94], N654, N651);
  xnor KeyGate_0_94(N727, keyIn_0_94, KeyWire_0[94]);
nor NOR2_253 (N731, N341, N659);
nand NAND2_254 (N732, N654, N261);
  nand NAND3_255 (KeyWire_0[95], N644, N654, N261);
  xor KeyGate_0_95(N733, keyIn_0_95, KeyWire_0[95]);
  nand NAND4_256 (KeyWire_0[96], N635, N644, N654, N261);
  xnor KeyGate_0_96(N734, keyIn_0_96, KeyWire_0[96]);
not NOT1_257 (N735, N662);
and AND2_258 (N736, N228, N665);
and AND2_259 (N737, N237, N662);
not NOT1_260 (N738, N670);
and AND2_261 (N739, N228, N673);
and AND2_262 (N740, N237, N670);
not NOT1_263 (N741, N678);
and AND2_264 (N742, N228, N682);
and AND2_265 (N743, N237, N678);
not NOT1_266 (N744, N687);
and AND2_267 (N745, N228, N692);
and AND2_268 (N746, N237, N687);
not NOT1_269 (N747, N697);
and AND2_270 (N748, N228, N700);
and AND2_271 (N749, N237, N697);
not NOT1_272 (N750, N705);
and AND2_273 (N751, N228, N708);
and AND2_274 (N752, N237, N705);
not NOT1_275 (N753, N713);
and AND2_276 (N754, N228, N717);
and AND2_277 (N755, N237, N713);
not NOT1_278 (N756, N722);
nor NOR2_279 (N757, N727, N261);
and AND2_280 (N758, N727, N261);
and AND2_281 (N759, N228, N727);
and AND2_282 (N760, N237, N722);
  nand NAND2_283 (KeyWire_0[97], N644, N722);
  xor KeyGate_0_97(KeyNOTWire_0[48], keyIn_0_97, KeyWire_0[97]);
  not KeyNOTGate_0_48(N761, KeyNOTWire_0[48]);
  nand NAND2_284 (KeyWire_0[98], N635, N713);
  xnor KeyGate_0_98(N762, keyIn_0_98, KeyWire_0[98]);
  nand NAND3_285 (KeyWire_0[99], N635, N644, N722);
  xnor KeyGate_0_99(KeyNOTWire_0[49], keyIn_0_99, KeyWire_0[99]);
  not KeyNOTGate_0_49(N763, KeyNOTWire_0[49]);
  nand NAND2_286 (KeyWire_0[100], N609, N687);
  xor KeyGate_0_100(N764, keyIn_0_100, KeyWire_0[100]);
  nand NAND2_287 (KeyWire_0[101], N600, N678);
  xnor KeyGate_0_101(KeyNOTWire_0[50], keyIn_0_101, KeyWire_0[101]);
  not KeyNOTGate_0_50(N765, KeyNOTWire_0[50]);
  nand NAND3_288 (KeyWire_0[102], N600, N609, N687);
  xor KeyGate_0_102(KeyNOTWire_0[51], keyIn_0_102, KeyWire_0[102]);
  not KeyNOTGate_0_51(N766, KeyNOTWire_0[51]);
buf BUFF1_289 (N767, N660);
buf BUFF1_290 (N768, N661);
nor NOR2_291 (N769, N736, N737);
nor NOR2_292 (N770, N739, N740);
nor NOR2_293 (N771, N742, N743);
nor NOR2_294 (N772, N745, N746);
  nand NAND4_295 (KeyWire_0[103], N750, N762, N763, N734);
  xor KeyGate_0_103(KeyNOTWire_0[52], keyIn_0_103, KeyWire_0[103]);
  not KeyNOTGate_0_52(N773, KeyNOTWire_0[52]);
nor NOR2_296 (N777, N748, N749);
  nand NAND3_297 (KeyWire_0[104], N753, N761, N733);
  xnor KeyGate_0_104(N778, keyIn_0_104, KeyWire_0[104]);
nor NOR2_298 (N781, N751, N752);
  nand NAND2_299 (KeyWire_0[105], N756, N732);
  xor KeyGate_0_105(N782, keyIn_0_105, KeyWire_0[105]);
nor NOR2_300 (N785, N754, N755);
nor NOR2_301 (N786, N757, N758);
nor NOR2_302 (N787, N759, N760);
nor NOR2_303 (N788, N700, N773);
  and AND2_304 (KeyWire_0[106], N700, N773);
  xnor KeyGate_0_106(N789, keyIn_0_106, KeyWire_0[106]);
nor NOR2_305 (N790, N708, N778);
  and AND2_306 (KeyWire_0[107], N708, N778);
  xor KeyGate_0_107(N791, keyIn_0_107, KeyWire_0[107]);
nor NOR2_307 (N792, N717, N782);
  and AND2_308 (KeyWire_0[108], N717, N782);
  xnor KeyGate_0_108(N793, keyIn_0_108, KeyWire_0[108]);
and AND2_309 (N794, N219, N786);
  nand NAND2_310 (KeyWire_0[109], N628, N773);
  xor KeyGate_0_109(N795, keyIn_0_109, KeyWire_0[109]);
  nand NAND2_311 (KeyWire_0[110], N795, N747);
  xnor KeyGate_0_110(N796, keyIn_0_110, KeyWire_0[110]);
nor NOR2_312 (N802, N788, N789);
nor NOR2_313 (N803, N790, N791);
nor NOR2_314 (N804, N792, N793);
nor NOR2_315 (N805, N340, N794);
nor NOR2_316 (N806, N692, N796);
  and AND2_317 (KeyWire_0[111], N692, N796);
  xnor KeyGate_0_111(KeyNOTWire_0[53], keyIn_0_111, KeyWire_0[111]);
  not KeyNOTGate_0_53(N807, KeyNOTWire_0[53]);
and AND2_318 (N808, N219, N802);
and AND2_319 (N809, N219, N803);
and AND2_320 (N810, N219, N804);
  nand NAND4_321 (KeyWire_0[112], N805, N787, N731, N529);
  xnor KeyGate_0_112(KeyNOTWire_0[54], keyIn_0_112, KeyWire_0[112]);
  not KeyNOTGate_0_54(N811, KeyNOTWire_0[54]);
  nand NAND2_322 (KeyWire_0[113], N619, N796);
  xnor KeyGate_0_113(N812, keyIn_0_113, KeyWire_0[113]);
  nand NAND3_323 (KeyWire_0[114], N609, N619, N796);
  xor KeyGate_0_114(KeyNOTWire_0[55], keyIn_0_114, KeyWire_0[114]);
  not KeyNOTGate_0_55(N813, KeyNOTWire_0[55]);
  nand NAND4_324 (KeyWire_0[115], N600, N609, N619, N796);
  xor KeyGate_0_115(N814, keyIn_0_115, KeyWire_0[115]);
  nand NAND4_325 (KeyWire_0[116], N738, N765, N766, N814);
  xnor KeyGate_0_116(KeyNOTWire_0[56], keyIn_0_116, KeyWire_0[116]);
  not KeyNOTGate_0_56(N815, KeyNOTWire_0[56]);
  nand NAND3_326 (KeyWire_0[117], N741, N764, N813);
  xor KeyGate_0_117(KeyNOTWire_0[57], keyIn_0_117, KeyWire_0[117]);
  not KeyNOTGate_0_57(N819, KeyNOTWire_0[57]);
  nand NAND2_327 (KeyWire_0[118], N744, N812);
  xor KeyGate_0_118(KeyNOTWire_0[58], keyIn_0_118, KeyWire_0[118]);
  not KeyNOTGate_0_58(N822, KeyNOTWire_0[58]);
nor NOR2_328 (N825, N806, N807);
nor NOR2_329 (N826, N335, N808);
nor NOR2_330 (N827, N336, N809);
nor NOR2_331 (N828, N338, N810);
not NOT1_332 (N829, N811);
nor NOR2_333 (N830, N665, N815);
and AND2_334 (N831, N665, N815);
nor NOR2_335 (N832, N673, N819);
  and AND2_336 (KeyWire_0[119], N673, N819);
  xnor KeyGate_0_119(N833, keyIn_0_119, KeyWire_0[119]);
nor NOR2_337 (N834, N682, N822);
  and AND2_338 (KeyWire_0[120], N682, N822);
  xor KeyGate_0_120(N835, keyIn_0_120, KeyWire_0[120]);
and AND2_339 (N836, N219, N825);
  nand NAND3_340 (KeyWire_0[121], N826, N777, N704);
  xor KeyGate_0_121(N837, keyIn_0_121, KeyWire_0[121]);
  nand NAND4_341 (KeyWire_0[122], N827, N781, N712, N527);
  xor KeyGate_0_122(KeyNOTWire_0[59], keyIn_0_122, KeyWire_0[122]);
  not KeyNOTGate_0_59(N838, KeyNOTWire_0[59]);
  nand NAND4_342 (KeyWire_0[123], N828, N785, N721, N528);
  xor KeyGate_0_123(KeyNOTWire_0[60], keyIn_0_123, KeyWire_0[123]);
  not KeyNOTGate_0_60(N839, KeyNOTWire_0[60]);
not NOT1_343 (N840, N829);
nand NAND2_344 (N841, N815, N593);
nor NOR2_345 (N842, N830, N831);
nor NOR2_346 (N843, N832, N833);
nor NOR2_347 (N844, N834, N835);
nor NOR2_348 (N845, N334, N836);
not NOT1_349 (N846, N837);
not NOT1_350 (N847, N838);
not NOT1_351 (N848, N839);
and AND2_352 (N849, N735, N841);
buf BUFF1_353 (N850, N840);
and AND2_354 (N851, N219, N842);
and AND2_355 (N852, N219, N843);
and AND2_356 (N853, N219, N844);
  nand NAND3_357 (KeyWire_0[124], N845, N772, N696);
  xnor KeyGate_0_124(KeyNOTWire_0[61], keyIn_0_124, KeyWire_0[124]);
  not KeyNOTGate_0_61(N854, KeyNOTWire_0[61]);
not NOT1_358 (N855, N846);
not NOT1_359 (N856, N847);
not NOT1_360 (N857, N848);
not NOT1_361 (N858, N849);
nor NOR2_362 (N859, N417, N851);
nor NOR2_363 (N860, N332, N852);
nor NOR2_364 (N861, N333, N853);
not NOT1_365 (N862, N854);
buf BUFF1_366 (N863, N855);
buf BUFF1_367 (N864, N856);
buf BUFF1_368 (N865, N857);
buf BUFF1_369 (N866, N858);
  nand NAND3_370 (KeyWire_0[125], N859, N769, N669);
  xnor KeyGate_0_125(N867, keyIn_0_125, KeyWire_0[125]);
  nand NAND3_371 (KeyWire_0[126], N860, N770, N677);
  xnor KeyGate_0_126(KeyNOTWire_0[62], keyIn_0_126, KeyWire_0[126]);
  not KeyNOTGate_0_62(N868, KeyNOTWire_0[62]);
  nand NAND3_372 (KeyWire_0[127], N861, N771, N686);
  xnor KeyGate_0_127(KeyNOTWire_0[63], keyIn_0_127, KeyWire_0[127]);
  not KeyNOTGate_0_63(N869, KeyNOTWire_0[63]);
not NOT1_373 (N870, N862);
not NOT1_374 (N871, N867);
not NOT1_375 (N872, N868);
not NOT1_376 (N873, N869);
buf BUFF1_377 (N874, N870);
not NOT1_378 (N875, N871);
not NOT1_379 (N876, N872);
not NOT1_380 (N877, N873);
buf BUFF1_381 (N878, N875);
buf BUFF1_382 (N879, N876);
buf BUFF1_383 (N880, N877);

endmodule
