`timescale 1ns / 1ps
// Verilog
// c880
// Ninputs 60
// Noutputs 26
// NtotalGates 383
// NAND4 13
// AND3 12
// NAND2 60
// NAND3 14
// AND2 105
// OR2 29
// NOT1 63
// NOR2 61
// BUFF1 26

module top (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
                  N865,N866,N874,N878,N879,N880,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
                  keyinput30, keyinput31,
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36,
        keyinput37, keyinput38, keyinput39, keyinput40, keyinput41,
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46,
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51,
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56,
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61,
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66,
        keyinput67, keyinput68, keyinput69, keyinput70, keyinput71,
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76,
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81,
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86,
        keyinput87, keyinput88, keyinput89, keyinput90, keyinput91,
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96,
        keyinput97, keyinput98, keyinput99, keyinput100, keyinput101,
        keyinput102, keyinput103, keyinput104, keyinput105, keyinput106,
        keyinput107, keyinput108, keyinput109, keyinput110, keyinput111,
        keyinput112, keyinput113, keyinput114, keyinput115, keyinput116,
        keyinput117, keyinput118, keyinput119, keyinput120, keyinput121,
        keyinput122, keyinput123, keyinput124, keyinput125, keyinput126,
        keyinput127, keyinput128, keyinput129, keyinput130, keyinput131,
        keyinput132, keyinput133, keyinput134, keyinput135, keyinput136,
        keyinput137, keyinput138, keyinput139, keyinput140, keyinput141,
        keyinput142, keyinput143, keyinput144, keyinput145, keyinput146,
                  keyinput147, keyinput148, keyinput149, keyinput150, keyinput151,
        keyinput152, keyinput153, keyinput154, keyinput155, keyinput156,
        keyinput157, keyinput158, keyinput159, keyinput160, keyinput161,
        keyinput162, keyinput163, keyinput164, keyinput165, keyinput166,
        keyinput167, keyinput168, keyinput169, keyinput170, keyinput171,
        keyinput172, keyinput173, keyinput174, keyinput175, keyinput176,
        keyinput177, keyinput178, keyinput179, keyinput180, keyinput181,
        keyinput182, keyinput183, keyinput184, keyinput185, keyinput186,
        keyinput187, keyinput188, keyinput189, keyinput190, keyinput191,
        keyinput192, keyinput193, keyinput194, keyinput195, keyinput196,
        keyinput197, keyinput198, keyinput199, keyinput200, keyinput201,
        keyinput202, keyinput203, keyinput204, keyinput205, keyinput206,
        keyinput207, keyinput208, keyinput209, keyinput210, keyinput211);

  input keyinput152, keyinput153, keyinput154, keyinput155, keyinput156;
  input keyinput157, keyinput158, keyinput159, keyinput160, keyinput161;
  input keyinput162, keyinput163, keyinput164, keyinput165, keyinput166;
  input keyinput167, keyinput168, keyinput169, keyinput170, keyinput171;
  input keyinput172, keyinput173, keyinput174, keyinput175, keyinput176;
  input keyinput177, keyinput178, keyinput179, keyinput180, keyinput181;
  input keyinput182, keyinput183, keyinput184, keyinput185, keyinput186;
  input keyinput187, keyinput188, keyinput189, keyinput190, keyinput191;
  input keyinput192, keyinput193, keyinput194, keyinput195, keyinput196;
  input keyinput197, keyinput198, keyinput199, keyinput200, keyinput201;
  input keyinput202, keyinput203, keyinput204, keyinput205, keyinput206;
  input keyinput207, keyinput208, keyinput209, keyinput210, keyinput211;


  input keyinput32, keyinput33, keyinput34, keyinput35, keyinput36;
  input keyinput37, keyinput38, keyinput39, keyinput40, keyinput41;
  input keyinput42, keyinput43, keyinput44, keyinput45, keyinput46;
  input keyinput47, keyinput48, keyinput49, keyinput50, keyinput51;
  input keyinput52, keyinput53, keyinput54, keyinput55, keyinput56;
  input keyinput57, keyinput58, keyinput59, keyinput60, keyinput61;
  input keyinput62, keyinput63, keyinput64, keyinput65, keyinput66;
  input keyinput67, keyinput68, keyinput69, keyinput70, keyinput71;
  input keyinput72, keyinput73, keyinput74, keyinput75, keyinput76;
  input keyinput77, keyinput78, keyinput79, keyinput80, keyinput81;
  input keyinput82, keyinput83, keyinput84, keyinput85, keyinput86;
  input keyinput87, keyinput88, keyinput89, keyinput90, keyinput91;
  input keyinput92, keyinput93, keyinput94, keyinput95, keyinput96;
  input keyinput97, keyinput98, keyinput99, keyinput100, keyinput101;
  input keyinput102, keyinput103, keyinput104, keyinput105, keyinput106;
  input keyinput107, keyinput108, keyinput109, keyinput110, keyinput111;
  input keyinput112, keyinput113, keyinput114, keyinput115, keyinput116;
  input keyinput117, keyinput118, keyinput119, keyinput120, keyinput121;
  input keyinput122, keyinput123, keyinput124, keyinput125, keyinput126;
  input keyinput127, keyinput128, keyinput129, keyinput130, keyinput131;
  input keyinput132, keyinput133, keyinput134, keyinput135, keyinput136;
  input keyinput137, keyinput138, keyinput139, keyinput140, keyinput141;
  input keyinput142, keyinput143, keyinput144, keyinput145, keyinput146;
  input keyinput147, keyinput148, keyinput149, keyinput150, keyinput151;

  wire KeyWire_0_1 , KeyWire_0_2, keyinput_Wire_1;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31;

  wire [0:31] keyinput_Wire_0;
  wire [0:16] KeyNOTWire_0;

input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;

output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;

wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877;

nand NAND4_1 (N269, N1, N8, N13, N17);
nand NAND4_2 (N270, N1, N26, N13, N17);
and AND3_3 (N273, N29, N36, N42);
and AND3_4 (N276, N1, N26, N51);
nand NAND4_5 (N279, N1, N8, N51, N17);
  nand NAND4_6 (keyinput_Wire_0[0], N1, N8, N13, N55);
  xnor keyGate_0_0(N280, keyinput0, keyinput_Wire_0[0]);
nand NAND4_7 (N284, N59, N42, N68, N72);
nand NAND2_8 (N285, N29, N68);
nand NAND3_9 (N286, N59, N68, N74);
  and AND3_10 (keyinput_Wire_0[1], N29, N75, N80);
  xor keyGate_0_1(N287, keyinput1, keyinput_Wire_0[1]);
and AND3_11 (N290, N29, N75, N42);
and AND3_12 (N291, N29, N36, N80);
and AND3_13 (N292, N29, N36, N42);
and AND3_14 (N293, N59, N75, N80);
and AND3_15 (N294, N59, N75, N42);
and AND3_16 (N295, N59, N36, N80);
and AND3_17 (N296, N59, N36, N42);
and AND2_18 (N297, N85, N86);
or OR2_19 (N298, N87, N88);
nand NAND2_20 (N301, N91, N96);
  or OR2_21 (keyinput_Wire_0[2], N91, N96);
  xnor keyGate_0_2(N302, keyinput2, keyinput_Wire_0[2]);
nand NAND2_22 (N303, N101, N106);
or OR2_23 (N304, N101, N106);
nand NAND2_24 (N305, N111, N116);
or OR2_25 (N306, N111, N116);
nand NAND2_26 (N307, N121, N126);
or OR2_27 (N308, N121, N126);
and AND2_28 (N309, N8, N138);
not NOT1_29 (N310, N268);
and AND2_30 (N316, N51, N138);
and AND2_31 (N317, N17, N138);
and AND2_32 (N318, N152, N138);
nand NAND2_33 (N319, N59, N156);
nor NOR2_34 (N322, N17, N42);
and AND2_35 (N323, N17, N42);
  nand NAND2_36 (keyinput_Wire_0[3], N159, N165);
  xnor keyGate_0_3(KeyNOTWire_0[0], keyinput3, keyinput_Wire_0[3]);
  not KeyNOTGate_0_0(N324, KeyNOTWire_0[0]);
or OR2_37 (N325, N159, N165);
nand NAND2_38 (N326, N171, N177);
or OR2_39 (N327, N171, N177);
nand NAND2_40 (N328, N183, N189);
or OR2_41 (N329, N183, N189);
  nand NAND2_42 (keyinput_Wire_0[4], N195, N201);
  xor keyGate_0_4(N330, keyinput4, keyinput_Wire_0[4]);
or OR2_43 (N331, N195, N201);
and AND2_44 (N332, N210, N91);
and AND2_45 (N333, N210, N96);
and AND2_46 (N334, N210, N101);
and AND2_47 (N335, N210, N106);
and AND2_48 (N336, N210, N111);
  and AND2_49 (keyinput_Wire_0[5], N255, N259);
  xor keyGate_0_5(KeyNOTWire_0[1], keyinput5, keyinput_Wire_0[5]);
  not KeyNOTGate_0_1(N337, KeyNOTWire_0[1]);
and AND2_50 (N338, N210, N116);
and AND2_51 (N339, N255, N260);
and AND2_52 (N340, N210, N121);
and AND2_53 (N341, N255, N267);
  not NOT1_54 (keyinput_Wire_0[6], N269);
  xnor keyGate_0_6(KeyNOTWire_0[2], keyinput6, keyinput_Wire_0[6]);
  not KeyNOTGate_0_2(N342, KeyNOTWire_0[2]);
  not NOT1_55 (keyinput_Wire_0[7], N273);
  xor keyGate_0_7(KeyNOTWire_0[3], keyinput7, keyinput_Wire_0[7]);
  not KeyNOTGate_0_3(N343, KeyNOTWire_0[3]);
or OR2_56 (N344, N270, N273);
not NOT1_57 (N345, N276);
not NOT1_58 (N346, N276);
not NOT1_59 (N347, N279);
nor NOR2_60 (N348, N280, N284);
or OR2_61 (N349, N280, N285);
or OR2_62 (N350, N280, N286);
not NOT1_63 (N351, N293);
not NOT1_64 (N352, N294);
not NOT1_65 (N353, N295);
not NOT1_66 (N354, N296);
nand NAND2_67 (N355, N89, N298);
and AND2_68 (N356, N90, N298);
nand NAND2_69 (N357, N301, N302);
nand NAND2_70 (N360, N303, N304);
nand NAND2_71 (N363, N305, N306);
  nand NAND2_72 (keyinput_Wire_0[8], N307, N308);
  xnor keyGate_0_8(KeyNOTWire_0[4], keyinput8, keyinput_Wire_0[8]);
  not KeyNOTGate_0_4(N366, KeyNOTWire_0[4]);
not NOT1_73 (N369, N310);
nor NOR2_74 (N375, N322, N323);
nand NAND2_75 (N376, N324, N325);
nand NAND2_76 (N379, N326, N327);
nand NAND2_77 (N382, N328, N329);
nand NAND2_78 (N385, N330, N331);
buf BUFF1_79 (N388, N290);
buf BUFF1_80 (N389, N291);
buf BUFF1_81 (N390, N292);
buf BUFF1_82 (N391, N297);
or OR2_83 (N392, N270, N343);
not NOT1_84 (N393, N345);
not NOT1_85 (N399, N346);
and AND2_86 (N400, N348, N73);
not NOT1_87 (N401, N349);
not NOT1_88 (N402, N350);
not NOT1_89 (N403, N355);
not NOT1_90 (N404, N357);
  not NOT1_91 (keyinput_Wire_0[9], N360);
  xor keyGate_0_9(N405, keyinput9, keyinput_Wire_0[9]);
  and AND2_92 (keyinput_Wire_0[10], N357, N360);
  xnor keyGate_0_10(KeyNOTWire_0[5], keyinput10, keyinput_Wire_0[10]);
  not KeyNOTGate_0_5(N406, KeyNOTWire_0[5]);
not NOT1_93 (N407, N363);
not NOT1_94 (N408, N366);
and AND2_95 (N409, N363, N366);
nand NAND2_96 (N410, N347, N352);
not NOT1_97 (N411, N376);
not NOT1_98 (N412, N379);
and AND2_99 (N413, N376, N379);
  not NOT1_100 (keyinput_Wire_0[11], N382);
  xnor keyGate_0_11(KeyNOTWire_0[6], keyinput11, keyinput_Wire_0[11]);
  not KeyNOTGate_0_6(N414, KeyNOTWire_0[6]);
  not NOT1_101 (keyinput_Wire_0[12], N385);
  xor keyGate_0_12(KeyNOTWire_0[7], keyinput12, keyinput_Wire_0[12]);
  not KeyNOTGate_0_7(N415, KeyNOTWire_0[7]);
and AND2_102 (N416, N382, N385);
and AND2_103 (N417, N210, N369);
buf BUFF1_104 (N418, N342);
buf BUFF1_105 (N419, N344);
buf BUFF1_106 (N420, N351);
buf BUFF1_107 (N421, N353);
buf BUFF1_108 (N422, N354);
buf BUFF1_109 (N423, N356);
not NOT1_110 (N424, N400);
and AND2_111 (N425, N404, N405);
and AND2_112 (N426, N407, N408);
  and AND3_113 (keyinput_Wire_0[13], N319, N393, N55);
  xnor keyGate_0_13(KeyNOTWire_0[8], keyinput13, keyinput_Wire_0[13]);
  not KeyNOTGate_0_8(N427, KeyNOTWire_0[8]);
and AND3_114 (N432, N393, N17, N287);
nand NAND3_115 (N437, N393, N287, N55);
nand NAND4_116 (N442, N375, N59, N156, N393);
nand NAND3_117 (N443, N393, N319, N17);
and AND2_118 (N444, N411, N412);
and AND2_119 (N445, N414, N415);
buf BUFF1_120 (N446, N392);
buf BUFF1_121 (N447, N399);
buf BUFF1_122 (N448, N401);
buf BUFF1_123 (N449, N402);
buf BUFF1_124 (N450, N403);
not NOT1_125 (N451, N424);
nor NOR2_126 (N460, N406, N425);
nor NOR2_127 (N463, N409, N426);
nand NAND2_128 (N466, N442, N410);
and AND2_129 (N475, N143, N427);
and AND2_130 (N476, N310, N432);
and AND2_131 (N477, N146, N427);
and AND2_132 (N478, N310, N432);
and AND2_133 (N479, N149, N427);
and AND2_134 (N480, N310, N432);
and AND2_135 (N481, N153, N427);
and AND2_136 (N482, N310, N432);
nand NAND2_137 (N483, N443, N1);
or OR2_138 (N488, N369, N437);
or OR2_139 (N489, N369, N437);
or OR2_140 (N490, N369, N437);
or OR2_141 (N491, N369, N437);
nor NOR2_142 (N492, N413, N444);
nor NOR2_143 (N495, N416, N445);
nand NAND2_144 (N498, N130, N460);
or OR2_145 (N499, N130, N460);
nand NAND2_146 (N500, N463, N135);
or OR2_147 (N501, N463, N135);
  and AND2_148 (keyinput_Wire_0[14], N91, N466);
  xnor keyGate_0_14(N502, keyinput14, keyinput_Wire_0[14]);
nor NOR2_149 (N503, N475, N476);
and AND2_150 (N504, N96, N466);
nor NOR2_151 (N505, N477, N478);
and AND2_152 (N506, N101, N466);
nor NOR2_153 (N507, N479, N480);
  and AND2_154 (keyinput_Wire_0[15], N106, N466);
  xnor keyGate_0_15(KeyNOTWire_0[9], keyinput15, keyinput_Wire_0[15]);
  not KeyNOTGate_0_9(N508, KeyNOTWire_0[9]);
nor NOR2_155 (N509, N481, N482);
and AND2_156 (N510, N143, N483);
and AND2_157 (N511, N111, N466);
and AND2_158 (N512, N146, N483);
and AND2_159 (N513, N116, N466);
  and AND2_160 (keyinput_Wire_0[16], N149, N483);
  xnor keyGate_0_16(KeyNOTWire_0[10], keyinput16, keyinput_Wire_0[16]);
  not KeyNOTGate_0_10(N514, KeyNOTWire_0[10]);
  and AND2_161 (keyinput_Wire_0[17], N121, N466);
  xnor keyGate_0_17(KeyNOTWire_0[11], keyinput17, keyinput_Wire_0[17]);
  not KeyNOTGate_0_11(N515, KeyNOTWire_0[11]);
and AND2_162 (N516, N153, N483);
and AND2_163 (N517, N126, N466);
nand NAND2_164 (N518, N130, N492);
or OR2_165 (N519, N130, N492);
nand NAND2_166 (N520, N495, N207);
or OR2_167 (N521, N495, N207);
and AND2_168 (N522, N451, N159);
and AND2_169 (N523, N451, N165);
and AND2_170 (N524, N451, N171);
and AND2_171 (N525, N451, N177);
and AND2_172 (N526, N451, N183);
nand NAND2_173 (N527, N451, N189);
nand NAND2_174 (N528, N451, N195);
nand NAND2_175 (N529, N451, N201);
nand NAND2_176 (N530, N498, N499);
nand NAND2_177 (N533, N500, N501);
nor NOR2_178 (N536, N309, N502);
nor NOR2_179 (N537, N316, N504);
nor NOR2_180 (N538, N317, N506);
nor NOR2_181 (N539, N318, N508);
nor NOR2_182 (N540, N510, N511);
nor NOR2_183 (N541, N512, N513);
  nor NOR2_184 (keyinput_Wire_0[18], N514, N515);
  xnor keyGate_0_18(KeyNOTWire_0[12], keyinput18, keyinput_Wire_0[18]);
  not KeyNOTGate_0_12(N542, KeyNOTWire_0[12]);
nor NOR2_185 (N543, N516, N517);
nand NAND2_186 (N544, N518, N519);
nand NAND2_187 (N547, N520, N521);
not NOT1_188 (N550, N530);
not NOT1_189 (N551, N533);
and AND2_190 (N552, N530, N533);
nand NAND2_191 (N553, N536, N503);
nand NAND2_192 (N557, N537, N505);
nand NAND2_193 (N561, N538, N507);
nand NAND2_194 (N565, N539, N509);
nand NAND2_195 (N569, N488, N540);
nand NAND2_196 (N573, N489, N541);
nand NAND2_197 (N577, N490, N542);
nand NAND2_198 (N581, N491, N543);
not NOT1_199 (N585, N544);
not NOT1_200 (N586, N547);
and AND2_201 (N587, N544, N547);
and AND2_202 (N588, N550, N551);
and AND2_203 (N589, N585, N586);
nand NAND2_204 (N590, N553, N159);
or OR2_205 (N593, N553, N159);
and AND2_206 (N596, N246, N553);
nand NAND2_207 (N597, N557, N165);
  or OR2_208 (keyinput_Wire_0[19], N557, N165);
  xnor keyGate_0_19(KeyNOTWire_0[13], keyinput19, keyinput_Wire_0[19]);
  not KeyNOTGate_0_13(N600, KeyNOTWire_0[13]);
and AND2_209 (N605, N246, N557);
nand NAND2_210 (N606, N561, N171);
or OR2_211 (N609, N561, N171);
and AND2_212 (N615, N246, N561);
nand NAND2_213 (N616, N565, N177);
or OR2_214 (N619, N565, N177);
and AND2_215 (N624, N246, N565);
nand NAND2_216 (N625, N569, N183);
or OR2_217 (N628, N569, N183);
and AND2_218 (N631, N246, N569);
nand NAND2_219 (N632, N573, N189);
or OR2_220 (N635, N573, N189);
and AND2_221 (N640, N246, N573);
nand NAND2_222 (N641, N577, N195);
or OR2_223 (N644, N577, N195);
and AND2_224 (N650, N246, N577);
nand NAND2_225 (N651, N581, N201);
or OR2_226 (N654, N581, N201);
  and AND2_227 (keyinput_Wire_0[20], N246, N581);
  xor keyGate_0_20(N659, keyinput20, keyinput_Wire_0[20]);
nor NOR2_228 (N660, N552, N588);
nor NOR2_229 (N661, N587, N589);
  not NOT1_230 (keyinput_Wire_0[21], N590);
  xnor keyGate_0_21(N662, keyinput21, keyinput_Wire_0[21]);
and AND2_231 (N665, N593, N590);
nor NOR2_232 (N669, N596, N522);
not NOT1_233 (N670, N597);
and AND2_234 (N673, N600, N597);
nor NOR2_235 (N677, N605, N523);
not NOT1_236 (N678, N606);
and AND2_237 (N682, N609, N606);
nor NOR2_238 (N686, N615, N524);
not NOT1_239 (N687, N616);
and AND2_240 (N692, N619, N616);
nor NOR2_241 (N696, N624, N525);
not NOT1_242 (N697, N625);
and AND2_243 (N700, N628, N625);
nor NOR2_244 (N704, N631, N526);
not NOT1_245 (N705, N632);
and AND2_246 (N708, N635, N632);
nor NOR2_247 (N712, N337, N640);
not NOT1_248 (N713, N641);
and AND2_249 (N717, N644, N641);
nor NOR2_250 (N721, N339, N650);
not NOT1_251 (N722, N651);
and AND2_252 (N727, N654, N651);
nor NOR2_253 (N731, N341, N659);
nand NAND2_254 (N732, N654, N261);
nand NAND3_255 (N733, N644, N654, N261);
nand NAND4_256 (N734, N635, N644, N654, N261);
not NOT1_257 (N735, N662);
and AND2_258 (N736, N228, N665);
  and AND2_259 (keyinput_Wire_0[22], N237, N662);
  xnor keyGate_0_22(KeyNOTWire_0[14], keyinput22, keyinput_Wire_0[22]);
  not KeyNOTGate_0_14(N737, KeyNOTWire_0[14]);
not NOT1_260 (N738, N670);
and AND2_261 (N739, N228, N673);
and AND2_262 (N740, N237, N670);
not NOT1_263 (N741, N678);
and AND2_264 (N742, N228, N682);
and AND2_265 (N743, N237, N678);
not NOT1_266 (N744, N687);
and AND2_267 (N745, N228, N692);
and AND2_268 (N746, N237, N687);
not NOT1_269 (N747, N697);
and AND2_270 (N748, N228, N700);
  and AND2_271 (keyinput_Wire_0[23], N237, N697);
  xnor keyGate_0_23(KeyNOTWire_0[15], keyinput23, keyinput_Wire_0[23]);
  not KeyNOTGate_0_15(N749, KeyNOTWire_0[15]);
not NOT1_272 (N750, N705);
and AND2_273 (N751, N228, N708);
  and AND2_274 (keyinput_Wire_0[24], N237, N705);
  xnor keyGate_0_24(N752, keyinput24, keyinput_Wire_0[24]);
not NOT1_275 (N753, N713);
and AND2_276 (N754, N228, N717);
and AND2_277 (N755, N237, N713);
not NOT1_278 (N756, N722);
nor NOR2_279 (N757, N727, N261);
  and AND2_280 (keyinput_Wire_0[25], N727, N261);
  xor keyGate_0_25(N758, keyinput25, keyinput_Wire_0[25]);
and AND2_281 (N759, N228, N727);
and AND2_282 (N760, N237, N722);
nand NAND2_283 (N761, N644, N722);
nand NAND2_284 (N762, N635, N713);
nand NAND3_285 (N763, N635, N644, N722);
nand NAND2_286 (N764, N609, N687);
nand NAND2_287 (N765, N600, N678);
nand NAND3_288 (N766, N600, N609, N687);
buf BUFF1_289 (N767, N660);
buf BUFF1_290 (N768, N661);
nor NOR2_291 (N769, N736, N737);
nor NOR2_292 (N770, N739, N740);
nor NOR2_293 (N771, N742, N743);
nor NOR2_294 (N772, N745, N746);
nand NAND4_295 (N773, N750, N762, N763, N734);
nor NOR2_296 (N777, N748, N749);
nand NAND3_297 (N778, N753, N761, N733);
nor NOR2_298 (N781, N751, N752);
nand NAND2_299 (N782, N756, N732);
  nor NOR2_300 (keyinput_Wire_0[26], N754, N755);
  xor keyGate_0_26(KeyNOTWire_0[16], keyinput26, keyinput_Wire_0[26]);
  not KeyNOTGate_0_16(N785, KeyNOTWire_0[16]);
nor NOR2_301 (N786, N757, N758);
nor NOR2_302 (N787, N759, N760);
nor NOR2_303 (N788, N700, N773);
and AND2_304 (N789, N700, N773);
nor NOR2_305 (N790, N708, N778);
and AND2_306 (N791, N708, N778);
nor NOR2_307 (N792, N717, N782);
and AND2_308 (N793, N717, N782);
and AND2_309 (N794, N219, N786);
nand NAND2_310 (N795, N628, N773);
nand NAND2_311 (N796, N795, N747);
nor NOR2_312 (N802, N788, N789);
  nor NOR2_313 (keyinput_Wire_0[27], N790, N791);
  xnor keyGate_0_27(N803, keyinput27, keyinput_Wire_0[27]);
nor NOR2_314 (N804, N792, N793);
  nor NOR2_315 (keyinput_Wire_0[28], N340, N794);
  xnor keyGate_0_28(N805, keyinput28, keyinput_Wire_0[28]);
nor NOR2_316 (N806, N692, N796);
and AND2_317 (N807, N692, N796);
and AND2_318 (N808, N219, N802);
and AND2_319 (N809, N219, N803);
and AND2_320 (N810, N219, N804);
nand NAND4_321 (N811, N805, N787, N731, N529);
nand NAND2_322 (N812, N619, N796);
nand NAND3_323 (N813, N609, N619, N796);
nand NAND4_324 (N814, N600, N609, N619, N796);
nand NAND4_325 (N815, N738, N765, N766, N814);
nand NAND3_326 (N819, N741, N764, N813);
nand NAND2_327 (N822, N744, N812);
nor NOR2_328 (N825, N806, N807);
nor NOR2_329 (N826, N335, N808);
nor NOR2_330 (N827, N336, N809);
nor NOR2_331 (N828, N338, N810);
not NOT1_332 (N829, N811);
nor NOR2_333 (N830, N665, N815);
and AND2_334 (N831, N665, N815);
nor NOR2_335 (N832, N673, N819);
and AND2_336 (N833, N673, N819);
nor NOR2_337 (N834, N682, N822);
and AND2_338 (N835, N682, N822);
and AND2_339 (N836, N219, N825);
nand NAND3_340 (N837, N826, N777, N704);
nand NAND4_341 (N838, N827, N781, N712, N527);
nand NAND4_342 (N839, N828, N785, N721, N528);
not NOT1_343 (N840, N829);
nand NAND2_344 (N841, N815, N593);
nor NOR2_345 (N842, N830, N831);
nor NOR2_346 (N843, N832, N833);
nor NOR2_347 (N844, N834, N835);
nor NOR2_348 (N845, N334, N836);
not NOT1_349 (N846, N837);
not NOT1_350 (N847, N838);
not NOT1_351 (N848, N839);
and AND2_352 (N849, N735, N841);
buf BUFF1_353 (N850, N840);
and AND2_354 (N851, N219, N842);
and AND2_355 (N852, N219, N843);
and AND2_356 (N853, N219, N844);
nand NAND3_357 (N854, N845, N772, N696);
not NOT1_358 (N855, N846);
not NOT1_359 (N856, N847);
not NOT1_360 (N857, N848);
not NOT1_361 (N858, N849);
  nor NOR2_362 (keyinput_Wire_0[29], N417, N851);
  xnor keyGate_0_29(N859, keyinput29, keyinput_Wire_0[29]);
nor NOR2_363 (N860, N332, N852);
nor NOR2_364 (N861, N333, N853);
not NOT1_365 (N862, N854);
buf BUFF1_366 (N863, N855);
buf BUFF1_367 (N864, N856);
  buf BUFF1_368 (keyinput_Wire_1, N857);
  xor keyGate_1_8(N865, KeyWire_0_2, keyinput_Wire_1);
buf BUFF1_369 (N866, N858);
nand NAND3_370 (N867, N859, N769, N669);
nand NAND3_371 (N868, N860, N770, N677);
nand NAND3_372 (N869, N861, N771, N686);
  not NOT1_373 (keyinput_Wire_0[30], N862);
  xor keyGate_0_30(N870, keyinput30, keyinput_Wire_0[30]);
  not NOT1_374 (keyinput_Wire_0[31], N867);
  xor keyGate_0_31(N871, keyinput31, keyinput_Wire_0[31]);
not NOT1_375 (N872, N868);
not NOT1_376 (N873, N869);
buf BUFF1_377 (N874, N870);
not NOT1_378 (N875, N871);
not NOT1_379 (N876, N872);
not NOT1_380 (N877, N873);
buf BUFF1_381 (N878, N875);
buf BUFF1_382 (N879, N876);
buf BUFF1_383 (N880, N877);

AntiSAT some_name( KeyWire_0_2, N68, N219, N42, N207, N51, N138, N259, N74, N55, N91, N268, N143, N255, N75, N152, N130, N146, N29, N1, N73, N201, N26, N17, N237, N149, N246, N88, N135, N183, N165, N171, N85, N106, N72, N159, N189, N101, N195, N59, N8, N36, N261, N86, N87, N80, N116, N156, N210, N121, N177, N228, N96, N267, N126, N260, N90, N89, N111, N153, N13, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151,
       keyinput152, keyinput153, keyinput154, keyinput155, keyinput156,
       keyinput157, keyinput158, keyinput159, keyinput160, keyinput161,
       keyinput162, keyinput163, keyinput164, keyinput165, keyinput166,
       keyinput167, keyinput168, keyinput169, keyinput170, keyinput171,
       keyinput172, keyinput173, keyinput174, keyinput175, keyinput176,
       keyinput177, keyinput178, keyinput179, keyinput180, keyinput181,
       keyinput182, keyinput183, keyinput184, keyinput185, keyinput186,
       keyinput187, keyinput188, keyinput189, keyinput190, keyinput191,
       keyinput192, keyinput193, keyinput194, keyinput195, keyinput196,
       keyinput197, keyinput198, keyinput199, keyinput200, keyinput201,
       keyinput202, keyinput203, keyinput204, keyinput205, keyinput206,
       keyinput207, keyinput208, keyinput209, keyinput210, keyinput211);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N68, N219, N42, N207, N51, N138, N259, N74, N55, N91, N268, N143, N255, N75, N152, N130, N146, N29, N1, N73, N201, N26, N17, N237, N149, N246, N88, N135, N183, N165, N171, N85, N106, N72, N159, N189, N101, N195, N59, N8, N36, N261, N86, N87, N80, N116, N156, N210, N121, N177, N228, N96, N267, N126, N260, N90, N89, N111, N153, N13, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151 ,
        keyinput152, keyinput153, keyinput154, keyinput155, keyinput156,
        keyinput157, keyinput158, keyinput159, keyinput160, keyinput161,
        keyinput162, keyinput163, keyinput164, keyinput165, keyinput166,
        keyinput167, keyinput168, keyinput169, keyinput170, keyinput171,
        keyinput172, keyinput173, keyinput174, keyinput175, keyinput176,
        keyinput177, keyinput178, keyinput179, keyinput180, keyinput181,
        keyinput182, keyinput183, keyinput184, keyinput185, keyinput186,
        keyinput187, keyinput188, keyinput189, keyinput190, keyinput191,
        keyinput192, keyinput193, keyinput194, keyinput195, keyinput196,
        keyinput197, keyinput198, keyinput199, keyinput200, keyinput201,
        keyinput202, keyinput203, keyinput204, keyinput205, keyinput206,
        keyinput207, keyinput208, keyinput209, keyinput210, keyinput211);

  input keyinput152, keyinput153, keyinput154, keyinput155, keyinput156;
  input keyinput157, keyinput158, keyinput159, keyinput160, keyinput161;
  input keyinput162, keyinput163, keyinput164, keyinput165, keyinput166;
  input keyinput167, keyinput168, keyinput169, keyinput170, keyinput171;
  input keyinput172, keyinput173, keyinput174, keyinput175, keyinput176;
  input keyinput177, keyinput178, keyinput179, keyinput180, keyinput181;
  input keyinput182, keyinput183, keyinput184, keyinput185, keyinput186;
  input keyinput187, keyinput188, keyinput189, keyinput190, keyinput191;
  input keyinput192, keyinput193, keyinput194, keyinput195, keyinput196;
  input keyinput197, keyinput198, keyinput199, keyinput200, keyinput201;
  input keyinput202, keyinput203, keyinput204, keyinput205, keyinput206;
  input keyinput207, keyinput208, keyinput209, keyinput210, keyinput211;

  wire [0:59] keyNTin_Wire_1;
  wire [0:30] KeyNOTWire_1;

  input N68, N219, N42, N207, N51, N138, N259, N74, N55, N91, N268, N143, N255, N75, N152, N130, N146, N29, N1, N73, N201, N26, N17, N237, N149, N246, N88, N135, N183, N165, N171, N85, N106, N72, N159, N189, N101, N195, N59, N8, N36, N261, N86, N87, N80, N116, N156, N210, N121, N177, N228, N96, N267, N126, N260, N90, N89, N111, N153, N13;
  input keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83, newWire_84, newWire_85, newWire_86, newWire_87, newWire_88, newWire_89, newWire_90, newWire_91, newWire_92, newWire_93, newWire_94, newWire_95, newWire_96, newWire_97, newWire_98, newWire_99, newWire_100, newWire_101, newWire_102, newWire_103, newWire_104, newWire_105, newWire_106, newWire_107, newWire_108, newWire_109, newWire_110, newWire_111, newWire_112, newWire_113, newWire_114, newWire_115, newWire_116, newWire_117, newWire_118, newWire_119, newWire_120, newWire_121 ;

  xor  KeyGate0 (keyNTin_Wire_1[0], N68, keyinput32);
  xnor keyNTinGate_1_0(newWire_0, keyinput152, keyNTin_Wire_1[0]);
  xor  KeyGate1 (newWire_1, N219, keyinput33);
  xor  KeyGate2 (keyNTin_Wire_1[1], N42, keyinput34);
  xnor keyNTinGate_1_1(newWire_2, keyinput153, keyNTin_Wire_1[1]);
  xnor KeyGate3 (keyNTin_Wire_1[2], N207, keyinput35);
  xor keyNTinGate_1_2(KeyNOTWire_1[0], keyinput154, keyNTin_Wire_1[2]);
  not KeyNOTGate_1_0(newWire_3, KeyNOTWire_1[0]);
  xnor KeyGate4 (newWire_4, N51, keyinput36);
  xor  KeyGate5 (keyNTin_Wire_1[3], N138, keyinput37);
  xor keyNTinGate_1_3(KeyNOTWire_1[1], keyinput155, keyNTin_Wire_1[3]);
  not KeyNOTGate_1_1(newWire_5, KeyNOTWire_1[1]);
  xnor KeyGate6 (newWire_6, N259, keyinput38);
  xor  KeyGate7 (keyNTin_Wire_1[4], N74, keyinput39);
  xor keyNTinGate_1_4(newWire_7, keyinput156, keyNTin_Wire_1[4]);
  xor  KeyGate8 (newWire_8, N55, keyinput40);
  xor  KeyGate9 (keyNTin_Wire_1[5], N91, keyinput41);
  xor keyNTinGate_1_5(KeyNOTWire_1[2], keyinput157, keyNTin_Wire_1[5]);
  not KeyNOTGate_1_2(newWire_9, KeyNOTWire_1[2]);
  xor  KeyGate10 (keyNTin_Wire_1[6], N268, keyinput42);
  xnor keyNTinGate_1_6(KeyNOTWire_1[3], keyinput158, keyNTin_Wire_1[6]);
  not KeyNOTGate_1_3(newWire_10, KeyNOTWire_1[3]);
  xor  KeyGate11 (newWire_11, N143, keyinput43);
  xnor KeyGate12 (newWire_12, N255, keyinput44);
  xor  KeyGate13 (keyNTin_Wire_1[7], N75, keyinput45);
  xor keyNTinGate_1_7(newWire_13, keyinput159, keyNTin_Wire_1[7]);
  xor  KeyGate14 (keyNTin_Wire_1[8], N152, keyinput46);
  xnor keyNTinGate_1_8(newWire_14, keyinput160, keyNTin_Wire_1[8]);
  xor  KeyGate15 (newWire_15, N130, keyinput47);
  xor  KeyGate16 (keyNTin_Wire_1[9], N146, keyinput48);
  xnor keyNTinGate_1_9(KeyNOTWire_1[4], keyinput161, keyNTin_Wire_1[9]);
  not KeyNOTGate_1_4(newWire_16, KeyNOTWire_1[4]);
  xor  KeyGate17 (newWire_17, N29, keyinput49);
  xnor KeyGate18 (newWire_18, N1, keyinput50);
  xnor KeyGate19 (newWire_19, N73, keyinput51);
  xnor KeyGate20 (keyNTin_Wire_1[10], N201, keyinput52);
  xor keyNTinGate_1_10(newWire_20, keyinput162, keyNTin_Wire_1[10]);
  xor  KeyGate21 (keyNTin_Wire_1[11], N26, keyinput53);
  xor keyNTinGate_1_11(newWire_21, keyinput163, keyNTin_Wire_1[11]);
  xor  KeyGate22 (newWire_22, N17, keyinput54);
  xnor KeyGate23 (keyNTin_Wire_1[12], N237, keyinput55);
  xnor keyNTinGate_1_12(KeyNOTWire_1[5], keyinput164, keyNTin_Wire_1[12]);
  not KeyNOTGate_1_5(newWire_23, KeyNOTWire_1[5]);
  xnor KeyGate24 (keyNTin_Wire_1[13], N149, keyinput56);
  xor keyNTinGate_1_13(KeyNOTWire_1[6], keyinput165, keyNTin_Wire_1[13]);
  not KeyNOTGate_1_6(newWire_24, KeyNOTWire_1[6]);
  xor  KeyGate25 (newWire_25, N246, keyinput57);
  xor  KeyGate26 (keyNTin_Wire_1[14], N88, keyinput58);
  xor keyNTinGate_1_14(newWire_26, keyinput166, keyNTin_Wire_1[14]);
  xnor KeyGate27 (keyNTin_Wire_1[15], N135, keyinput59);
  xor keyNTinGate_1_15(KeyNOTWire_1[7], keyinput167, keyNTin_Wire_1[15]);
  not KeyNOTGate_1_7(newWire_27, KeyNOTWire_1[7]);
  xnor KeyGate28 (keyNTin_Wire_1[16], N183, keyinput60);
  xnor keyNTinGate_1_16(newWire_28, keyinput168, keyNTin_Wire_1[16]);
  xnor KeyGate29 (newWire_29, N165, keyinput61);
  xnor KeyGate30 (keyNTin_Wire_1[17], N171, keyinput62);
  xor keyNTinGate_1_17(newWire_30, keyinput169, keyNTin_Wire_1[17]);
  xor  KeyGate31 (keyNTin_Wire_1[18], N85, keyinput63);
  xor keyNTinGate_1_18(KeyNOTWire_1[8], keyinput170, keyNTin_Wire_1[18]);
  not KeyNOTGate_1_8(newWire_31, KeyNOTWire_1[8]);
  xnor KeyGate32 (newWire_32, N106, keyinput64);
  xnor KeyGate33 (newWire_33, N72, keyinput65);
  xor  KeyGate34 (keyNTin_Wire_1[19], N159, keyinput66);
  xnor keyNTinGate_1_19(KeyNOTWire_1[9], keyinput171, keyNTin_Wire_1[19]);
  not KeyNOTGate_1_9(newWire_34, KeyNOTWire_1[9]);
  xor  KeyGate35 (keyNTin_Wire_1[20], N189, keyinput67);
  xnor keyNTinGate_1_20(newWire_35, keyinput172, keyNTin_Wire_1[20]);
  xor  KeyGate36 (newWire_36, N101, keyinput68);
  xor  KeyGate37 (keyNTin_Wire_1[21], N195, keyinput69);
  xor keyNTinGate_1_21(newWire_37, keyinput173, keyNTin_Wire_1[21]);
  xnor KeyGate38 (newWire_38, N59, keyinput70);
  xor  KeyGate39 (keyNTin_Wire_1[22], N8, keyinput71);
  xnor keyNTinGate_1_22(newWire_39, keyinput174, keyNTin_Wire_1[22]);
  xnor KeyGate40 (keyNTin_Wire_1[23], N36, keyinput72);
  xor keyNTinGate_1_23(KeyNOTWire_1[10], keyinput175, keyNTin_Wire_1[23]);
  not KeyNOTGate_1_10(newWire_40, KeyNOTWire_1[10]);
  xor  KeyGate41 (newWire_41, N261, keyinput73);
  xnor KeyGate42 (newWire_42, N86, keyinput74);
  xnor KeyGate43 (newWire_43, N87, keyinput75);
  xor  KeyGate44 (keyNTin_Wire_1[24], N80, keyinput76);
  xnor keyNTinGate_1_24(KeyNOTWire_1[11], keyinput176, keyNTin_Wire_1[24]);
  not KeyNOTGate_1_11(newWire_44, KeyNOTWire_1[11]);
  xor  KeyGate45 (keyNTin_Wire_1[25], N116, keyinput77);
  xnor keyNTinGate_1_25(KeyNOTWire_1[12], keyinput177, keyNTin_Wire_1[25]);
  not KeyNOTGate_1_12(newWire_45, KeyNOTWire_1[12]);
  xnor KeyGate46 (newWire_46, N156, keyinput78);
  xor  KeyGate47 (newWire_47, N210, keyinput79);
  xor  KeyGate48 (keyNTin_Wire_1[26], N121, keyinput80);
  xnor keyNTinGate_1_26(KeyNOTWire_1[13], keyinput178, keyNTin_Wire_1[26]);
  not KeyNOTGate_1_13(newWire_48, KeyNOTWire_1[13]);
  xor  KeyGate49 (keyNTin_Wire_1[27], N177, keyinput81);
  xor keyNTinGate_1_27(KeyNOTWire_1[14], keyinput179, keyNTin_Wire_1[27]);
  not KeyNOTGate_1_14(newWire_49, KeyNOTWire_1[14]);
  xnor KeyGate50 (newWire_50, N228, keyinput82);
  xor  KeyGate51 (keyNTin_Wire_1[28], N96, keyinput83);
  xnor keyNTinGate_1_28(KeyNOTWire_1[15], keyinput180, keyNTin_Wire_1[28]);
  not KeyNOTGate_1_15(newWire_51, KeyNOTWire_1[15]);
  xor  KeyGate52 (newWire_52, N267, keyinput84);
  xor  KeyGate53 (keyNTin_Wire_1[29], N126, keyinput85);
  xor keyNTinGate_1_29(newWire_53, keyinput181, keyNTin_Wire_1[29]);
  xnor KeyGate54 (keyNTin_Wire_1[30], N260, keyinput86);
  xor keyNTinGate_1_30(newWire_54, keyinput182, keyNTin_Wire_1[30]);
  xnor KeyGate55 (keyNTin_Wire_1[31], N90, keyinput87);
  xor keyNTinGate_1_31(newWire_55, keyinput183, keyNTin_Wire_1[31]);
  xnor KeyGate56 (newWire_56, N89, keyinput88);
  xor  KeyGate57 (newWire_57, N111, keyinput89);
  xnor KeyGate58 (newWire_58, N153, keyinput90);
  xnor KeyGate59 (newWire_59, N13, keyinput91);
  xnor KeyGate60 (newWire_60, N68, keyinput92);
  xor  KeyGate61 (newWire_61, N219, keyinput93);
  xnor KeyGate62 (keyNTin_Wire_1[32], N42, keyinput94);
  xor keyNTinGate_1_32(KeyNOTWire_1[16], keyinput184, keyNTin_Wire_1[32]);
  not KeyNOTGate_1_16(newWire_62, KeyNOTWire_1[16]);
  xnor KeyGate63 (keyNTin_Wire_1[33], N207, keyinput95);
  xor keyNTinGate_1_33(newWire_63, keyinput185, keyNTin_Wire_1[33]);
  xnor KeyGate64 (newWire_64, N51, keyinput96);
  xnor KeyGate65 (keyNTin_Wire_1[34], N138, keyinput97);
  xor keyNTinGate_1_34(newWire_65, keyinput186, keyNTin_Wire_1[34]);
  xor  KeyGate66 (keyNTin_Wire_1[35], N259, keyinput98);
  xnor keyNTinGate_1_35(KeyNOTWire_1[17], keyinput187, keyNTin_Wire_1[35]);
  not KeyNOTGate_1_17(newWire_66, KeyNOTWire_1[17]);
  xor  KeyGate67 (keyNTin_Wire_1[36], N74, keyinput99);
  xnor keyNTinGate_1_36(newWire_67, keyinput188, keyNTin_Wire_1[36]);
  xnor KeyGate68 (newWire_68, N55, keyinput100);
  xor  KeyGate69 (keyNTin_Wire_1[37], N91, keyinput101);
  xnor keyNTinGate_1_37(newWire_69, keyinput189, keyNTin_Wire_1[37]);
  xor  KeyGate70 (keyNTin_Wire_1[38], N268, keyinput102);
  xor keyNTinGate_1_38(newWire_70, keyinput190, keyNTin_Wire_1[38]);
  xnor KeyGate71 (newWire_71, N143, keyinput103);
  xor  KeyGate72 (keyNTin_Wire_1[39], N255, keyinput104);
  xnor keyNTinGate_1_39(KeyNOTWire_1[18], keyinput191, keyNTin_Wire_1[39]);
  not KeyNOTGate_1_18(newWire_72, KeyNOTWire_1[18]);
  xnor KeyGate73 (newWire_73, N75, keyinput105);
  xor  KeyGate74 (newWire_74, N152, keyinput106);
  xnor KeyGate75 (keyNTin_Wire_1[40], N130, keyinput107);
  xor keyNTinGate_1_40(newWire_75, keyinput192, keyNTin_Wire_1[40]);
  xnor KeyGate76 (newWire_76, N146, keyinput108);
  xnor KeyGate77 (keyNTin_Wire_1[41], N29, keyinput109);
  xnor keyNTinGate_1_41(KeyNOTWire_1[19], keyinput193, keyNTin_Wire_1[41]);
  not KeyNOTGate_1_19(newWire_77, KeyNOTWire_1[19]);
  xnor KeyGate78 (keyNTin_Wire_1[42], N1, keyinput110);
  xnor keyNTinGate_1_42(newWire_78, keyinput194, keyNTin_Wire_1[42]);
  xnor KeyGate79 (keyNTin_Wire_1[43], N73, keyinput111);
  xor keyNTinGate_1_43(newWire_79, keyinput195, keyNTin_Wire_1[43]);
  xor  KeyGate80 (newWire_80, N201, keyinput112);
  xnor KeyGate81 (keyNTin_Wire_1[44], N26, keyinput113);
  xnor keyNTinGate_1_44(KeyNOTWire_1[20], keyinput196, keyNTin_Wire_1[44]);
  not KeyNOTGate_1_20(newWire_81, KeyNOTWire_1[20]);
  xor  KeyGate82 (keyNTin_Wire_1[45], N17, keyinput114);
  xor keyNTinGate_1_45(KeyNOTWire_1[21], keyinput197, keyNTin_Wire_1[45]);
  not KeyNOTGate_1_21(newWire_82, KeyNOTWire_1[21]);
  xnor KeyGate83 (newWire_83, N237, keyinput115);
  xor  KeyGate84 (newWire_84, N149, keyinput116);
  xor  KeyGate85 (newWire_85, N246, keyinput117);
  xnor KeyGate86 (newWire_86, N88, keyinput118);
  xnor KeyGate87 (keyNTin_Wire_1[46], N135, keyinput119);
  xnor keyNTinGate_1_46(KeyNOTWire_1[22], keyinput198, keyNTin_Wire_1[46]);
  not KeyNOTGate_1_22(newWire_87, KeyNOTWire_1[22]);
  xor  KeyGate88 (newWire_88, N183, keyinput120);
  xnor KeyGate89 (keyNTin_Wire_1[47], N165, keyinput121);
  xnor keyNTinGate_1_47(KeyNOTWire_1[23], keyinput199, keyNTin_Wire_1[47]);
  not KeyNOTGate_1_23(newWire_89, KeyNOTWire_1[23]);
  xor  KeyGate90 (keyNTin_Wire_1[48], N171, keyinput122);
  xor keyNTinGate_1_48(newWire_90, keyinput200, keyNTin_Wire_1[48]);
  xnor KeyGate91 (keyNTin_Wire_1[49], N85, keyinput123);
  xor keyNTinGate_1_49(KeyNOTWire_1[24], keyinput201, keyNTin_Wire_1[49]);
  not KeyNOTGate_1_24(newWire_91, KeyNOTWire_1[24]);
  xor  KeyGate92 (newWire_92, N106, keyinput124);
  xnor KeyGate93 (keyNTin_Wire_1[50], N72, keyinput125);
  xor keyNTinGate_1_50(KeyNOTWire_1[25], keyinput202, keyNTin_Wire_1[50]);
  not KeyNOTGate_1_25(newWire_93, KeyNOTWire_1[25]);
  xnor KeyGate94 (newWire_94, N159, keyinput126);
  xnor KeyGate95 (keyNTin_Wire_1[51], N189, keyinput127);
  xnor keyNTinGate_1_51(KeyNOTWire_1[26], keyinput203, keyNTin_Wire_1[51]);
  not KeyNOTGate_1_26(newWire_95, KeyNOTWire_1[26]);
  xnor KeyGate96 (keyNTin_Wire_1[52], N101, keyinput128);
  xor keyNTinGate_1_52(newWire_96, keyinput204, keyNTin_Wire_1[52]);
  xor  KeyGate97 (keyNTin_Wire_1[53], N195, keyinput129);
  xnor keyNTinGate_1_53(KeyNOTWire_1[27], keyinput205, keyNTin_Wire_1[53]);
  not KeyNOTGate_1_27(newWire_97, KeyNOTWire_1[27]);
  xnor KeyGate98 (keyNTin_Wire_1[54], N59, keyinput130);
  xnor keyNTinGate_1_54(KeyNOTWire_1[28], keyinput206, keyNTin_Wire_1[54]);
  not KeyNOTGate_1_28(newWire_98, KeyNOTWire_1[28]);
  xnor KeyGate99 (newWire_99, N8, keyinput131);
  xor  KeyGate100 (newWire_100, N36, keyinput132);
  xnor KeyGate101 (newWire_101, N261, keyinput133);
  xor  KeyGate102 (newWire_102, N86, keyinput134);
  xnor KeyGate103 (newWire_103, N87, keyinput135);
  xor  KeyGate104 (newWire_104, N80, keyinput136);
  xnor KeyGate105 (newWire_105, N116, keyinput137);
  xor  KeyGate106 (keyNTin_Wire_1[55], N156, keyinput138);
  xnor keyNTinGate_1_55(KeyNOTWire_1[29], keyinput207, keyNTin_Wire_1[55]);
  not KeyNOTGate_1_29(newWire_106, KeyNOTWire_1[29]);
  xnor KeyGate107 (keyNTin_Wire_1[56], N210, keyinput139);
  xnor keyNTinGate_1_56(newWire_107, keyinput208, keyNTin_Wire_1[56]);
  xor  KeyGate108 (newWire_108, N121, keyinput140);
  xor  KeyGate109 (newWire_109, N177, keyinput141);
  xor  KeyGate110 (keyNTin_Wire_1[57], N228, keyinput142);
  xor keyNTinGate_1_57(newWire_110, keyinput209, keyNTin_Wire_1[57]);
  xnor KeyGate111 (newWire_111, N96, keyinput143);
  xor  KeyGate112 (newWire_112, N267, keyinput144);
  xnor KeyGate113 (newWire_113, N126, keyinput145);
  xnor KeyGate114 (newWire_114, N260, keyinput146);
  xor  KeyGate115 (keyNTin_Wire_1[58], N90, keyinput147);
  xnor keyNTinGate_1_58(newWire_115, keyinput210, keyNTin_Wire_1[58]);
  xnor KeyGate116 (keyNTin_Wire_1[59], N89, keyinput148);
  xnor keyNTinGate_1_59(KeyNOTWire_1[30], keyinput211, keyNTin_Wire_1[59]);
  not KeyNOTGate_1_30(newWire_116, KeyNOTWire_1[30]);
  xnor KeyGate117 (newWire_117, N111, keyinput149);
  xnor KeyGate118 (newWire_118, N153, keyinput150);
  xor  KeyGate119 (newWire_119, N13, keyinput151);
  and some_function (newWire_120, newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59 );
  nand compl_function (newWire_121, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83, newWire_84, newWire_85, newWire_86, newWire_87, newWire_88, newWire_89, newWire_90, newWire_91, newWire_92, newWire_93, newWire_94, newWire_95, newWire_96, newWire_97, newWire_98, newWire_99, newWire_100, newWire_101, newWire_102, newWire_103, newWire_104, newWire_105, newWire_106, newWire_107, newWire_108, newWire_109, newWire_110, newWire_111, newWire_112, newWire_113, newWire_114, newWire_115, newWire_116, newWire_117, newWire_118, newWire_119);
  and finalAND (KeyWire_0_2, newWire_120, newWire_121);

endmodule /* AntiSAT */
