// Benchmark "C432_locked" written by ABC on Wed Sep  6 17:13:42 2017

module top ( 
    G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat,
    G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat, G56gat,
    G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, G82gat, G86gat,
    G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, G108gat, G112gat,
    G115gat, keyinput0_G223gat, keyinput1_G223gat, keyinput2_G223gat,
    keyinput3_G223gat, keyinput0_G329gat, keyinput1_G329gat,
    keyinput2_G329gat, keyinput3_G329gat, keyinput0_G370gat,
    keyinput1_G370gat, keyinput2_G370gat, keyinput3_G370gat,
    keyinput0_G421gat, keyinput1_G421gat, keyinput2_G421gat,
    keyinput3_G421gat, keyinput0_G430gat, keyinput1_G430gat,
    keyinput2_G430gat, keyinput3_G430gat, keyinput0_G431gat,
    keyinput1_G431gat, keyinput2_G431gat, keyinput3_G431gat,
    keyinput0_G432gat, keyinput1_G432gat, keyinput2_G432gat,
    keyinput3_G432gat,
    G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat  );
  input  G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat,
    G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat,
    G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, G82gat,
    G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, G108gat,
    G112gat, G115gat, keyinput0_G223gat, keyinput1_G223gat,
    keyinput2_G223gat, keyinput3_G223gat, keyinput0_G329gat,
    keyinput1_G329gat, keyinput2_G329gat, keyinput3_G329gat,
    keyinput0_G370gat, keyinput1_G370gat, keyinput2_G370gat,
    keyinput3_G370gat, keyinput0_G421gat, keyinput1_G421gat,
    keyinput2_G421gat, keyinput3_G421gat, keyinput0_G430gat,
    keyinput1_G430gat, keyinput2_G430gat, keyinput3_G430gat,
    keyinput0_G431gat, keyinput1_G431gat, keyinput2_G431gat,
    keyinput3_G431gat, keyinput0_G432gat, keyinput1_G432gat,
    keyinput2_G432gat, keyinput3_G432gat;
  output G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat;
  wire n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
    n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
    n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
    n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
    n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
    n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
    n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
    n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
    n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
    n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
    n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
    n943, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
    n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
    n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
    n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
    n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
    n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
    n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
    n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
    n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
    n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
    n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
    n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
    n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
    n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
    n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
    n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
    n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
    n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
    n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
    n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
    n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
    n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
    n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
    n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
    n1313, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
    n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
    n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
    n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
    n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
    n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
    n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
    n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
    n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
    n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
    n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
    n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
    n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
    n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
    n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
    n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
    n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
    n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
    n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
    n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
    n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
    n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
    n1824, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
    n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
    n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
    n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
    n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
    n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
    n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
    n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
    n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
    n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
    n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
    n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
    n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
    n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
    n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
    n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
    n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
    n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
    n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
    n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
    n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
    n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
    n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
    n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
    n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
    n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
    n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
    n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
    n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
    n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
    n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
    n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
    n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
    n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
    n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
    n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
    n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
    n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
    n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
    n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
    n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
    n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
    n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
    n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
    n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
    n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
    n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
    n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
    n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
    n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
    n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
    n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
    n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
    n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
    n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
    n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
    n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
    n2445, n2446, n2447, n2448, n2449, n2450;
  assign n72 = ~G102gat & G108gat;
  assign n73 = ~G112gat & n72;
  assign n74 = ~G115gat & n73;
  assign n75 = G105gat & ~n74;
  assign n76 = ~G99gat & ~n75;
  assign n77 = ~G115gat & n72;
  assign n78 = ~G105gat & ~n73;
  assign n79 = ~n77 & ~n78;
  assign n80 = G99gat & ~n79;
  assign n81 = ~n76 & ~n80;
  assign n82 = ~keyinput0_G223gat & ~n81;
  assign n83 = keyinput0_G223gat & ~n75;
  assign n84 = ~n82 & ~n83;
  assign n85 = ~keyinput1_G223gat & ~n84;
  assign n86 = ~G108gat & ~G112gat;
  assign n87 = G112gat & ~n72;
  assign n88 = ~n86 & ~n87;
  assign n89 = G99gat & ~n88;
  assign n90 = ~keyinput0_G223gat & n89;
  assign n91 = G105gat & n74;
  assign n92 = ~G99gat & ~n91;
  assign n93 = G112gat & G115gat;
  assign n94 = n72 & ~n93;
  assign n95 = G105gat & ~n94;
  assign n96 = ~n78 & ~n95;
  assign n97 = G99gat & ~n96;
  assign n98 = ~n92 & ~n97;
  assign n99 = ~G89gat & ~n98;
  assign n100 = ~G105gat & ~n72;
  assign n101 = ~G112gat & ~G115gat;
  assign n102 = G102gat & ~n101;
  assign n103 = G108gat & ~n102;
  assign n104 = G105gat & ~n103;
  assign n105 = ~n100 & ~n104;
  assign n106 = ~G99gat & ~n105;
  assign n107 = ~G105gat & n89;
  assign n108 = ~n106 & ~n107;
  assign n109 = G89gat & ~n108;
  assign n110 = G102gat & n93;
  assign n111 = G108gat & ~n110;
  assign n112 = G105gat & ~n111;
  assign n113 = G89gat & G99gat;
  assign n114 = n112 & n113;
  assign n115 = ~n109 & ~n114;
  assign n116 = ~n99 & n115;
  assign n117 = keyinput0_G223gat & ~n116;
  assign n118 = ~n90 & ~n117;
  assign n119 = keyinput1_G223gat & ~n118;
  assign n120 = ~n85 & ~n119;
  assign n121 = ~keyinput2_G223gat & ~n120;
  assign n122 = G115gat & n72;
  assign n123 = ~G105gat & ~n122;
  assign n124 = G108gat & ~G115gat;
  assign n125 = G102gat & G112gat;
  assign n126 = n124 & ~n125;
  assign n127 = G105gat & n126;
  assign n128 = ~n123 & ~n127;
  assign n129 = ~G99gat & ~n128;
  assign n130 = G108gat & ~G112gat;
  assign n131 = G112gat & n72;
  assign n132 = ~n130 & ~n131;
  assign n133 = G115gat & ~n132;
  assign n134 = G99gat & ~n133;
  assign n135 = G105gat & ~n124;
  assign n136 = n134 & ~n135;
  assign n137 = ~n129 & ~n136;
  assign n138 = ~keyinput0_G223gat & ~n137;
  assign n139 = keyinput0_G223gat & ~n128;
  assign n140 = ~n138 & ~n139;
  assign n141 = ~keyinput1_G223gat & ~n140;
  assign n142 = G95gat & ~n113;
  assign n143 = ~n88 & ~n142;
  assign n144 = ~keyinput0_G223gat & n143;
  assign n145 = G99gat & ~n73;
  assign n146 = ~G89gat & ~n145;
  assign n147 = ~G99gat & ~n72;
  assign n148 = ~n130 & ~n147;
  assign n149 = G89gat & ~n148;
  assign n150 = ~n146 & ~n149;
  assign n151 = keyinput0_G223gat & ~n150;
  assign n152 = ~n144 & ~n151;
  assign n153 = keyinput1_G223gat & ~n152;
  assign n154 = ~n141 & ~n153;
  assign n155 = keyinput2_G223gat & ~n154;
  assign n156 = ~n121 & ~n155;
  assign n157 = ~keyinput3_G223gat & ~n156;
  assign n158 = G105gat & n113;
  assign n159 = G95gat & ~n158;
  assign n160 = ~n111 & ~n159;
  assign n161 = keyinput0_G223gat & n160;
  assign n162 = ~n90 & ~n161;
  assign n163 = ~keyinput1_G223gat & ~n162;
  assign n164 = ~keyinput0_G223gat & ~n112;
  assign n165 = keyinput0_G223gat & ~n111;
  assign n166 = ~n164 & ~n165;
  assign n167 = keyinput1_G223gat & ~n166;
  assign n168 = ~n163 & ~n167;
  assign n169 = ~keyinput2_G223gat & ~n168;
  assign n170 = G108gat & ~keyinput0_G223gat;
  assign n171 = ~G11gat & G17gat;
  assign n172 = ~G37gat & G43gat;
  assign n173 = ~G89gat & G95gat;
  assign n174 = ~G76gat & G82gat;
  assign n175 = ~n173 & ~n174;
  assign n176 = ~n72 & n175;
  assign n177 = ~G63gat & G69gat;
  assign n178 = ~G50gat & G56gat;
  assign n179 = ~n177 & ~n178;
  assign n180 = n176 & n179;
  assign n181 = ~n172 & n180;
  assign n182 = ~G24gat & G30gat;
  assign n183 = n181 & ~n182;
  assign n184 = ~G1gat & G4gat;
  assign n185 = n183 & ~n184;
  assign n186 = ~n171 & n185;
  assign n187 = keyinput0_G223gat & ~n186;
  assign n188 = ~n170 & ~n187;
  assign n189 = keyinput1_G223gat & ~n188;
  assign n190 = keyinput0_G223gat & ~n124;
  assign n191 = ~keyinput1_G223gat & ~n190;
  assign n192 = ~n170 & n191;
  assign n193 = ~n189 & ~n192;
  assign n194 = keyinput2_G223gat & ~n193;
  assign n195 = ~n169 & ~n194;
  assign n196 = keyinput3_G223gat & ~n195;
  assign G223gat = n157 | n196;
  assign n198 = ~keyinput3_G329gat & ~n79;
  assign n199 = keyinput3_G329gat & n160;
  assign n200 = ~n198 & ~n199;
  assign n201 = ~keyinput2_G329gat & ~n200;
  assign n202 = G89gat & ~n72;
  assign n203 = ~G89gat & ~G99gat;
  assign n204 = ~G102gat & ~G112gat;
  assign n205 = G108gat & n204;
  assign n206 = ~n203 & ~n205;
  assign n207 = ~n202 & n206;
  assign n208 = ~keyinput3_G329gat & ~n207;
  assign n209 = keyinput3_G329gat & ~n202;
  assign n210 = ~n208 & ~n209;
  assign n211 = keyinput2_G329gat & ~n210;
  assign n212 = ~n201 & ~n211;
  assign n213 = ~keyinput1_G329gat & ~n212;
  assign n214 = ~G89gat & G102gat;
  assign n215 = G105gat & ~G115gat;
  assign n216 = ~G99gat & ~n215;
  assign n217 = ~G112gat & ~n216;
  assign n218 = G99gat & n215;
  assign n219 = ~n217 & ~n218;
  assign n220 = ~n214 & ~n219;
  assign n221 = G89gat & ~G102gat;
  assign n222 = ~n220 & ~n221;
  assign n223 = G108gat & ~n222;
  assign n224 = ~keyinput3_G329gat & ~n223;
  assign n225 = keyinput3_G329gat & ~n112;
  assign n226 = ~n224 & ~n225;
  assign n227 = ~keyinput2_G329gat & ~n226;
  assign n228 = ~keyinput3_G329gat & n126;
  assign n229 = ~G108gat & keyinput3_G329gat;
  assign n230 = ~n228 & ~n229;
  assign n231 = keyinput2_G329gat & ~n230;
  assign n232 = ~n227 & ~n231;
  assign n233 = keyinput1_G329gat & ~n232;
  assign n234 = ~n213 & ~n233;
  assign n235 = ~keyinput0_G329gat & ~n234;
  assign n236 = G37gat & n179;
  assign n237 = n175 & n236;
  assign n238 = ~keyinput3_G329gat & ~n237;
  assign n239 = keyinput2_G329gat & ~n238;
  assign n240 = keyinput3_G329gat & n175;
  assign n241 = ~n239 & ~n240;
  assign n242 = ~n72 & ~n241;
  assign n243 = ~G99gat & ~G105gat;
  assign n244 = G89gat & ~n243;
  assign n245 = ~n103 & n244;
  assign n246 = ~keyinput3_G329gat & ~n245;
  assign n247 = ~keyinput2_G329gat & n246;
  assign n248 = ~n242 & ~n247;
  assign n249 = ~keyinput1_G329gat & n248;
  assign n250 = ~keyinput3_G329gat & n219;
  assign n251 = n72 & ~n250;
  assign n252 = ~keyinput2_G329gat & ~n251;
  assign n253 = G108gat & ~n125;
  assign n254 = ~keyinput3_G329gat & n253;
  assign n255 = G95gat & ~G99gat;
  assign n256 = ~G108gat & n255;
  assign n257 = ~G99gat & n173;
  assign n258 = G112gat & ~n257;
  assign n259 = ~G102gat & ~n258;
  assign n260 = ~G112gat & ~n173;
  assign n261 = ~n255 & ~n260;
  assign n262 = G102gat & ~n261;
  assign n263 = ~n259 & ~n262;
  assign n264 = G108gat & ~n263;
  assign n265 = ~n256 & ~n264;
  assign n266 = ~G82gat & ~n265;
  assign n267 = ~n205 & ~n257;
  assign n268 = G86gat & n267;
  assign n269 = ~G76gat & ~n268;
  assign n270 = ~n72 & ~n173;
  assign n271 = n267 & ~n270;
  assign n272 = ~G86gat & ~n271;
  assign n273 = G86gat & ~n265;
  assign n274 = ~n272 & ~n273;
  assign n275 = G76gat & ~n274;
  assign n276 = ~n269 & ~n275;
  assign n277 = G82gat & ~n276;
  assign n278 = ~n266 & ~n277;
  assign n279 = ~G69gat & ~n278;
  assign n280 = ~G76gat & ~G86gat;
  assign n281 = G82gat & n280;
  assign n282 = n267 & ~n281;
  assign n283 = G73gat & n282;
  assign n284 = ~G63gat & ~n283;
  assign n285 = ~n176 & n282;
  assign n286 = ~G73gat & ~n285;
  assign n287 = G73gat & ~n278;
  assign n288 = ~n286 & ~n287;
  assign n289 = G63gat & ~n288;
  assign n290 = ~n284 & ~n289;
  assign n291 = G69gat & ~n290;
  assign n292 = ~n279 & ~n291;
  assign n293 = ~G56gat & ~n292;
  assign n294 = ~G63gat & ~G73gat;
  assign n295 = G69gat & n294;
  assign n296 = n282 & ~n295;
  assign n297 = G60gat & n296;
  assign n298 = ~G50gat & ~n297;
  assign n299 = ~n177 & ~n285;
  assign n300 = G69gat & n284;
  assign n301 = ~n299 & ~n300;
  assign n302 = ~G60gat & ~n301;
  assign n303 = G60gat & ~n292;
  assign n304 = ~n302 & ~n303;
  assign n305 = G50gat & ~n304;
  assign n306 = ~n298 & ~n305;
  assign n307 = G56gat & ~n306;
  assign n308 = ~n293 & ~n307;
  assign n309 = ~G43gat & ~n308;
  assign n310 = ~G50gat & ~G60gat;
  assign n311 = G56gat & n310;
  assign n312 = n296 & ~n311;
  assign n313 = G47gat & n312;
  assign n314 = ~G37gat & ~n313;
  assign n315 = ~n178 & n301;
  assign n316 = n178 & n297;
  assign n317 = ~n315 & ~n316;
  assign n318 = ~G47gat & n317;
  assign n319 = G47gat & ~n308;
  assign n320 = ~n318 & ~n319;
  assign n321 = G37gat & ~n320;
  assign n322 = ~n314 & ~n321;
  assign n323 = G43gat & ~n322;
  assign n324 = ~n309 & ~n323;
  assign n325 = ~G30gat & ~n324;
  assign n326 = ~G37gat & ~G47gat;
  assign n327 = G43gat & n326;
  assign n328 = n312 & ~n327;
  assign n329 = G34gat & n328;
  assign n330 = ~G24gat & ~n329;
  assign n331 = ~n172 & ~n317;
  assign n332 = n172 & n313;
  assign n333 = ~n331 & ~n332;
  assign n334 = ~G34gat & n333;
  assign n335 = G34gat & ~n324;
  assign n336 = ~n334 & ~n335;
  assign n337 = G24gat & ~n336;
  assign n338 = ~n330 & ~n337;
  assign n339 = G30gat & ~n338;
  assign n340 = ~n325 & ~n339;
  assign n341 = ~G17gat & ~n340;
  assign n342 = ~G24gat & ~G34gat;
  assign n343 = G30gat & n342;
  assign n344 = n328 & ~n343;
  assign n345 = G21gat & n344;
  assign n346 = ~G11gat & ~n345;
  assign n347 = ~n182 & ~n333;
  assign n348 = n182 & n329;
  assign n349 = ~n347 & ~n348;
  assign n350 = ~G21gat & n349;
  assign n351 = G21gat & ~n340;
  assign n352 = ~n350 & ~n351;
  assign n353 = G11gat & ~n352;
  assign n354 = ~n346 & ~n353;
  assign n355 = G17gat & ~n354;
  assign n356 = ~n341 & ~n355;
  assign n357 = ~G4gat & ~n356;
  assign n358 = ~G11gat & ~G21gat;
  assign n359 = G17gat & n358;
  assign n360 = G8gat & n344;
  assign n361 = ~n359 & n360;
  assign n362 = ~G1gat & ~n361;
  assign n363 = ~G8gat & n349;
  assign n364 = G8gat & ~n340;
  assign n365 = ~n363 & ~n364;
  assign n366 = ~G17gat & ~n365;
  assign n367 = G21gat & ~n365;
  assign n368 = ~n350 & ~n367;
  assign n369 = G11gat & ~n368;
  assign n370 = ~n346 & ~n369;
  assign n371 = G17gat & ~n370;
  assign n372 = ~n366 & ~n371;
  assign n373 = G1gat & ~n372;
  assign n374 = ~n362 & ~n373;
  assign n375 = G4gat & ~n374;
  assign n376 = ~n357 & ~n375;
  assign n377 = keyinput3_G329gat & ~n376;
  assign n378 = ~n254 & ~n377;
  assign n379 = keyinput2_G329gat & ~n378;
  assign n380 = ~n252 & ~n379;
  assign n381 = keyinput1_G329gat & ~n380;
  assign n382 = ~n249 & ~n381;
  assign n383 = keyinput0_G329gat & ~n382;
  assign G329gat = n235 | n383;
  assign n385 = ~keyinput0_G370gat & ~n73;
  assign n386 = keyinput0_G370gat & n104;
  assign n387 = ~n385 & ~n386;
  assign n388 = ~keyinput1_G370gat & ~n387;
  assign n389 = ~G105gat & ~keyinput0_G370gat;
  assign n390 = n74 & ~n389;
  assign n391 = keyinput1_G370gat & ~n390;
  assign n392 = ~n388 & ~n391;
  assign n393 = ~keyinput2_G370gat & ~n392;
  assign n394 = ~G95gat & n130;
  assign n395 = G95gat & ~n150;
  assign n396 = ~n394 & ~n395;
  assign n397 = ~keyinput0_G370gat & ~n396;
  assign n398 = keyinput0_G370gat & ~n180;
  assign n399 = ~n397 & ~n398;
  assign n400 = ~keyinput1_G370gat & ~n399;
  assign n401 = keyinput0_G370gat & n72;
  assign n402 = ~keyinput0_G370gat & ~n132;
  assign n403 = ~n401 & ~n402;
  assign n404 = keyinput1_G370gat & ~n403;
  assign n405 = ~n400 & ~n404;
  assign n406 = keyinput2_G370gat & ~n405;
  assign n407 = ~n393 & ~n406;
  assign n408 = ~keyinput3_G370gat & ~n407;
  assign n409 = ~keyinput0_G370gat & n114;
  assign n410 = keyinput0_G370gat & ~n176;
  assign n411 = ~n409 & ~n410;
  assign n412 = ~keyinput1_G370gat & ~n411;
  assign n413 = ~keyinput0_G370gat & n112;
  assign n414 = ~n401 & ~n413;
  assign n415 = keyinput1_G370gat & n414;
  assign n416 = ~n412 & ~n415;
  assign n417 = ~keyinput2_G370gat & ~n416;
  assign n418 = ~keyinput0_G370gat & ~n202;
  assign n419 = ~n401 & ~n418;
  assign n420 = ~keyinput1_G370gat & ~n419;
  assign n421 = ~G108gat & ~keyinput0_G370gat;
  assign n422 = ~G95gat & n124;
  assign n423 = ~G89gat & ~n81;
  assign n424 = G89gat & ~n137;
  assign n425 = ~n423 & ~n424;
  assign n426 = G95gat & ~n425;
  assign n427 = ~n422 & ~n426;
  assign n428 = ~G82gat & ~n427;
  assign n429 = ~G89gat & n243;
  assign n430 = G95gat & n429;
  assign n431 = ~n74 & ~n430;
  assign n432 = G92gat & n431;
  assign n433 = ~G86gat & ~n432;
  assign n434 = G115gat & n73;
  assign n435 = ~n257 & n434;
  assign n436 = n75 & n257;
  assign n437 = ~n435 & ~n436;
  assign n438 = ~G92gat & n437;
  assign n439 = ~n77 & ~n173;
  assign n440 = n81 & n173;
  assign n441 = ~n439 & ~n440;
  assign n442 = G92gat & n441;
  assign n443 = ~n438 & ~n442;
  assign n444 = G86gat & ~n443;
  assign n445 = ~n433 & ~n444;
  assign n446 = ~G76gat & ~n445;
  assign n447 = n122 & ~n173;
  assign n448 = ~n440 & ~n447;
  assign n449 = ~G92gat & n448;
  assign n450 = ~G95gat & n126;
  assign n451 = G99gat & n126;
  assign n452 = ~n129 & ~n451;
  assign n453 = G89gat & ~n452;
  assign n454 = ~n423 & ~n453;
  assign n455 = G95gat & ~n454;
  assign n456 = ~n450 & ~n455;
  assign n457 = G92gat & ~n456;
  assign n458 = ~n449 & ~n457;
  assign n459 = ~G86gat & ~n458;
  assign n460 = ~G95gat & ~n133;
  assign n461 = ~n129 & ~n134;
  assign n462 = G89gat & ~n461;
  assign n463 = ~n423 & ~n462;
  assign n464 = G95gat & ~n463;
  assign n465 = ~n460 & ~n464;
  assign n466 = ~G92gat & ~n465;
  assign n467 = G92gat & ~n427;
  assign n468 = ~n466 & ~n467;
  assign n469 = G86gat & ~n468;
  assign n470 = ~n459 & ~n469;
  assign n471 = G76gat & ~n470;
  assign n472 = ~n446 & ~n471;
  assign n473 = G82gat & ~n472;
  assign n474 = ~n428 & ~n473;
  assign n475 = ~G69gat & ~n474;
  assign n476 = ~G86gat & ~G92gat;
  assign n477 = n174 & n476;
  assign n478 = n431 & ~n477;
  assign n479 = G79gat & n478;
  assign n480 = ~G73gat & ~n479;
  assign n481 = ~n281 & ~n437;
  assign n482 = n281 & n432;
  assign n483 = ~n481 & ~n482;
  assign n484 = ~G79gat & n483;
  assign n485 = ~n174 & n441;
  assign n486 = G82gat & n446;
  assign n487 = ~n485 & ~n486;
  assign n488 = G79gat & ~n487;
  assign n489 = ~n484 & ~n488;
  assign n490 = G73gat & ~n489;
  assign n491 = ~n480 & ~n490;
  assign n492 = ~G63gat & ~n491;
  assign n493 = ~n174 & n448;
  assign n494 = ~n486 & ~n493;
  assign n495 = ~G79gat & ~n494;
  assign n496 = ~G82gat & ~n456;
  assign n497 = G86gat & ~n456;
  assign n498 = ~n459 & ~n497;
  assign n499 = G76gat & ~n498;
  assign n500 = ~n446 & ~n499;
  assign n501 = G82gat & ~n500;
  assign n502 = ~n496 & ~n501;
  assign n503 = G79gat & ~n502;
  assign n504 = ~n495 & ~n503;
  assign n505 = ~G73gat & ~n504;
  assign n506 = ~G82gat & ~n465;
  assign n507 = G86gat & ~n465;
  assign n508 = ~n459 & ~n507;
  assign n509 = G76gat & ~n508;
  assign n510 = ~n446 & ~n509;
  assign n511 = G82gat & ~n510;
  assign n512 = ~n506 & ~n511;
  assign n513 = ~G79gat & ~n512;
  assign n514 = G79gat & ~n474;
  assign n515 = ~n513 & ~n514;
  assign n516 = G73gat & ~n515;
  assign n517 = ~n505 & ~n516;
  assign n518 = G63gat & ~n517;
  assign n519 = ~n492 & ~n518;
  assign n520 = G69gat & ~n519;
  assign n521 = ~n475 & ~n520;
  assign n522 = ~G56gat & ~n521;
  assign n523 = ~G73gat & ~G79gat;
  assign n524 = n177 & n523;
  assign n525 = n478 & ~n524;
  assign n526 = G66gat & n525;
  assign n527 = ~G60gat & ~n526;
  assign n528 = ~n295 & ~n483;
  assign n529 = n295 & n479;
  assign n530 = ~n528 & ~n529;
  assign n531 = ~G66gat & n530;
  assign n532 = ~n177 & ~n487;
  assign n533 = G69gat & n492;
  assign n534 = ~n532 & ~n533;
  assign n535 = G66gat & ~n534;
  assign n536 = ~n531 & ~n535;
  assign n537 = G60gat & ~n536;
  assign n538 = ~n527 & ~n537;
  assign n539 = ~G50gat & ~n538;
  assign n540 = ~n177 & ~n494;
  assign n541 = ~n533 & ~n540;
  assign n542 = ~G66gat & ~n541;
  assign n543 = ~G69gat & ~n502;
  assign n544 = G73gat & ~n502;
  assign n545 = ~n505 & ~n544;
  assign n546 = G63gat & ~n545;
  assign n547 = ~n492 & ~n546;
  assign n548 = G69gat & ~n547;
  assign n549 = ~n543 & ~n548;
  assign n550 = G66gat & ~n549;
  assign n551 = ~n542 & ~n550;
  assign n552 = ~G60gat & ~n551;
  assign n553 = ~G69gat & ~n512;
  assign n554 = G73gat & ~n512;
  assign n555 = ~n505 & ~n554;
  assign n556 = G63gat & ~n555;
  assign n557 = ~n492 & ~n556;
  assign n558 = G69gat & ~n557;
  assign n559 = ~n553 & ~n558;
  assign n560 = ~G66gat & ~n559;
  assign n561 = G66gat & ~n521;
  assign n562 = ~n560 & ~n561;
  assign n563 = G60gat & ~n562;
  assign n564 = ~n552 & ~n563;
  assign n565 = G50gat & ~n564;
  assign n566 = ~n539 & ~n565;
  assign n567 = G56gat & ~n566;
  assign n568 = ~n522 & ~n567;
  assign n569 = ~G43gat & ~n568;
  assign n570 = G56gat & ~G66gat;
  assign n571 = n310 & n570;
  assign n572 = n525 & ~n571;
  assign n573 = G53gat & n572;
  assign n574 = ~G47gat & ~n573;
  assign n575 = ~n311 & ~n530;
  assign n576 = n311 & n526;
  assign n577 = ~n575 & ~n576;
  assign n578 = ~G53gat & n577;
  assign n579 = ~n178 & ~n534;
  assign n580 = G56gat & n539;
  assign n581 = ~n579 & ~n580;
  assign n582 = G53gat & ~n581;
  assign n583 = ~n578 & ~n582;
  assign n584 = G47gat & ~n583;
  assign n585 = ~n574 & ~n584;
  assign n586 = ~G37gat & ~n585;
  assign n587 = ~n178 & ~n541;
  assign n588 = ~n580 & ~n587;
  assign n589 = ~G53gat & ~n588;
  assign n590 = ~G56gat & ~n549;
  assign n591 = G60gat & ~n549;
  assign n592 = ~n552 & ~n591;
  assign n593 = G50gat & ~n592;
  assign n594 = ~n539 & ~n593;
  assign n595 = G56gat & ~n594;
  assign n596 = ~n590 & ~n595;
  assign n597 = G53gat & ~n596;
  assign n598 = ~n589 & ~n597;
  assign n599 = ~G47gat & ~n598;
  assign n600 = ~G56gat & ~n559;
  assign n601 = G60gat & ~n559;
  assign n602 = ~n552 & ~n601;
  assign n603 = G50gat & ~n602;
  assign n604 = ~n539 & ~n603;
  assign n605 = G56gat & ~n604;
  assign n606 = ~n600 & ~n605;
  assign n607 = ~G53gat & ~n606;
  assign n608 = G53gat & ~n568;
  assign n609 = ~n607 & ~n608;
  assign n610 = G47gat & ~n609;
  assign n611 = ~n599 & ~n610;
  assign n612 = G37gat & ~n611;
  assign n613 = ~n586 & ~n612;
  assign n614 = G43gat & ~n613;
  assign n615 = ~n569 & ~n614;
  assign n616 = ~G30gat & ~n615;
  assign n617 = ~G47gat & ~G53gat;
  assign n618 = n172 & n617;
  assign n619 = n572 & ~n618;
  assign n620 = G40gat & n619;
  assign n621 = ~G34gat & ~n620;
  assign n622 = ~n327 & ~n577;
  assign n623 = n327 & n573;
  assign n624 = ~n622 & ~n623;
  assign n625 = ~G40gat & n624;
  assign n626 = ~n172 & ~n581;
  assign n627 = G43gat & n586;
  assign n628 = ~n626 & ~n627;
  assign n629 = G40gat & ~n628;
  assign n630 = ~n625 & ~n629;
  assign n631 = G34gat & ~n630;
  assign n632 = ~n621 & ~n631;
  assign n633 = ~G24gat & ~n632;
  assign n634 = ~n172 & ~n588;
  assign n635 = ~n627 & ~n634;
  assign n636 = ~G40gat & ~n635;
  assign n637 = ~G43gat & ~n596;
  assign n638 = G47gat & ~n596;
  assign n639 = ~n599 & ~n638;
  assign n640 = G37gat & ~n639;
  assign n641 = ~n586 & ~n640;
  assign n642 = G43gat & ~n641;
  assign n643 = ~n637 & ~n642;
  assign n644 = G40gat & ~n643;
  assign n645 = ~n636 & ~n644;
  assign n646 = ~G34gat & ~n645;
  assign n647 = ~G43gat & ~n606;
  assign n648 = G47gat & ~n606;
  assign n649 = ~n599 & ~n648;
  assign n650 = G37gat & ~n649;
  assign n651 = ~n586 & ~n650;
  assign n652 = G43gat & ~n651;
  assign n653 = ~n647 & ~n652;
  assign n654 = ~G40gat & ~n653;
  assign n655 = G40gat & ~n615;
  assign n656 = ~n654 & ~n655;
  assign n657 = G34gat & ~n656;
  assign n658 = ~n646 & ~n657;
  assign n659 = G24gat & ~n658;
  assign n660 = ~n633 & ~n659;
  assign n661 = G30gat & ~n660;
  assign n662 = ~n616 & ~n661;
  assign n663 = ~G17gat & ~n662;
  assign n664 = ~G34gat & ~G40gat;
  assign n665 = n182 & n664;
  assign n666 = n619 & ~n665;
  assign n667 = G27gat & n666;
  assign n668 = ~G21gat & ~n667;
  assign n669 = ~n343 & ~n624;
  assign n670 = n343 & n620;
  assign n671 = ~n669 & ~n670;
  assign n672 = ~G27gat & n671;
  assign n673 = ~n182 & ~n628;
  assign n674 = G30gat & n633;
  assign n675 = ~n673 & ~n674;
  assign n676 = G27gat & ~n675;
  assign n677 = ~n672 & ~n676;
  assign n678 = G21gat & ~n677;
  assign n679 = ~n668 & ~n678;
  assign n680 = ~G11gat & ~n679;
  assign n681 = ~n182 & ~n635;
  assign n682 = ~n674 & ~n681;
  assign n683 = ~G27gat & ~n682;
  assign n684 = ~G30gat & ~n643;
  assign n685 = G34gat & ~n643;
  assign n686 = ~n646 & ~n685;
  assign n687 = G24gat & ~n686;
  assign n688 = ~n633 & ~n687;
  assign n689 = G30gat & ~n688;
  assign n690 = ~n684 & ~n689;
  assign n691 = G27gat & ~n690;
  assign n692 = ~n683 & ~n691;
  assign n693 = ~G21gat & ~n692;
  assign n694 = ~G30gat & ~n653;
  assign n695 = G34gat & ~n653;
  assign n696 = ~n646 & ~n695;
  assign n697 = G24gat & ~n696;
  assign n698 = ~n633 & ~n697;
  assign n699 = G30gat & ~n698;
  assign n700 = ~n694 & ~n699;
  assign n701 = ~G27gat & ~n700;
  assign n702 = G27gat & ~n662;
  assign n703 = ~n701 & ~n702;
  assign n704 = G21gat & ~n703;
  assign n705 = ~n693 & ~n704;
  assign n706 = G11gat & ~n705;
  assign n707 = ~n680 & ~n706;
  assign n708 = G17gat & ~n707;
  assign n709 = ~n663 & ~n708;
  assign n710 = ~G4gat & ~n709;
  assign n711 = ~G14gat & ~n682;
  assign n712 = G14gat & ~n690;
  assign n713 = ~n711 & ~n712;
  assign n714 = ~G8gat & ~n713;
  assign n715 = ~G14gat & ~n700;
  assign n716 = G14gat & ~n662;
  assign n717 = ~n715 & ~n716;
  assign n718 = G8gat & ~n717;
  assign n719 = ~n714 & ~n718;
  assign n720 = ~G17gat & ~n719;
  assign n721 = G14gat & ~n692;
  assign n722 = ~n711 & ~n721;
  assign n723 = ~G21gat & ~n722;
  assign n724 = G21gat & ~n713;
  assign n725 = ~n723 & ~n724;
  assign n726 = ~G8gat & ~n725;
  assign n727 = G14gat & ~n703;
  assign n728 = ~n715 & ~n727;
  assign n729 = G21gat & ~n728;
  assign n730 = ~n693 & ~n729;
  assign n731 = G8gat & ~n730;
  assign n732 = ~n726 & ~n731;
  assign n733 = G11gat & ~n732;
  assign n734 = ~n680 & ~n733;
  assign n735 = G17gat & ~n734;
  assign n736 = ~n720 & ~n735;
  assign n737 = G1gat & ~n736;
  assign n738 = G14gat & n666;
  assign n739 = ~G8gat & ~n738;
  assign n740 = ~G14gat & n671;
  assign n741 = G14gat & ~n675;
  assign n742 = ~n740 & ~n741;
  assign n743 = G8gat & ~n742;
  assign n744 = ~n739 & ~n743;
  assign n745 = ~n171 & ~n744;
  assign n746 = G14gat & ~n677;
  assign n747 = ~n740 & ~n746;
  assign n748 = G21gat & ~n747;
  assign n749 = ~n668 & ~n748;
  assign n750 = G8gat & ~n749;
  assign n751 = ~G21gat & ~G27gat;
  assign n752 = n738 & ~n751;
  assign n753 = ~G8gat & ~n752;
  assign n754 = ~n750 & ~n753;
  assign n755 = n171 & ~n754;
  assign n756 = ~n745 & ~n755;
  assign n757 = ~G1gat & ~n756;
  assign n758 = ~n737 & ~n757;
  assign n759 = G4gat & ~n758;
  assign n760 = ~n710 & ~n759;
  assign n761 = keyinput0_G370gat & ~n760;
  assign n762 = ~n421 & ~n761;
  assign n763 = keyinput1_G370gat & ~n762;
  assign n764 = ~n420 & ~n763;
  assign n765 = keyinput2_G370gat & ~n764;
  assign n766 = ~n417 & ~n765;
  assign n767 = keyinput3_G370gat & ~n766;
  assign G370gat = n408 | n767;
  assign n769 = ~keyinput3_G421gat & ~n81;
  assign n770 = keyinput3_G421gat & n89;
  assign n771 = ~n769 & ~n770;
  assign n772 = ~keyinput2_G421gat & ~n771;
  assign n773 = ~keyinput3_G421gat & ~n137;
  assign n774 = ~G108gat & keyinput3_G421gat;
  assign n775 = ~n773 & ~n774;
  assign n776 = keyinput2_G421gat & ~n775;
  assign n777 = ~n772 & ~n776;
  assign n778 = ~keyinput1_G421gat & ~n777;
  assign n779 = ~keyinput3_G421gat & n89;
  assign n780 = keyinput3_G421gat & ~n112;
  assign n781 = ~n779 & ~n780;
  assign n782 = ~keyinput2_G421gat & ~n781;
  assign n783 = ~keyinput3_G421gat & ~n143;
  assign n784 = ~n774 & ~n783;
  assign n785 = keyinput2_G421gat & n784;
  assign n786 = ~n782 & ~n785;
  assign n787 = keyinput1_G421gat & ~n786;
  assign n788 = ~n778 & ~n787;
  assign n789 = ~keyinput0_G421gat & ~n788;
  assign n790 = ~keyinput3_G421gat & ~n75;
  assign n791 = keyinput3_G421gat & n160;
  assign n792 = ~n790 & ~n791;
  assign n793 = ~keyinput2_G421gat & ~n792;
  assign n794 = ~keyinput3_G421gat & ~n128;
  assign n795 = keyinput3_G421gat & n124;
  assign n796 = ~n794 & ~n795;
  assign n797 = keyinput2_G421gat & ~n796;
  assign n798 = ~n793 & ~n797;
  assign n799 = ~keyinput1_G421gat & ~n798;
  assign n800 = ~keyinput3_G421gat & ~n116;
  assign n801 = keyinput3_G421gat & ~n111;
  assign n802 = ~n800 & ~n801;
  assign n803 = ~keyinput2_G421gat & ~n802;
  assign n804 = ~keyinput3_G421gat & ~n150;
  assign n805 = ~G69gat & ~G82gat;
  assign n806 = ~G56gat & ~G108gat;
  assign n807 = n805 & n806;
  assign n808 = ~G43gat & ~G95gat;
  assign n809 = ~G17gat & ~G30gat;
  assign n810 = n808 & n809;
  assign n811 = n807 & n810;
  assign n812 = ~G4gat & ~n811;
  assign n813 = ~G14gat & ~n183;
  assign n814 = G76gat & ~n476;
  assign n815 = G82gat & ~n814;
  assign n816 = G63gat & ~n523;
  assign n817 = G69gat & ~n816;
  assign n818 = ~n815 & ~n817;
  assign n819 = G95gat & ~n244;
  assign n820 = ~G60gat & ~G66gat;
  assign n821 = G50gat & ~n820;
  assign n822 = G56gat & ~n821;
  assign n823 = G37gat & ~n617;
  assign n824 = G43gat & ~n823;
  assign n825 = G24gat & ~n664;
  assign n826 = G30gat & ~n825;
  assign n827 = ~n824 & ~n826;
  assign n828 = ~n822 & n827;
  assign n829 = ~n819 & n828;
  assign n830 = n818 & n829;
  assign n831 = ~n126 & n830;
  assign n832 = ~n122 & n831;
  assign n833 = G14gat & ~n832;
  assign n834 = ~n813 & ~n833;
  assign n835 = ~G8gat & ~n834;
  assign n836 = G76gat & G86gat;
  assign n837 = G82gat & ~n836;
  assign n838 = G63gat & G73gat;
  assign n839 = G69gat & ~n838;
  assign n840 = G50gat & G60gat;
  assign n841 = G56gat & ~n840;
  assign n842 = G37gat & G47gat;
  assign n843 = G43gat & ~n842;
  assign n844 = G24gat & G34gat;
  assign n845 = G30gat & ~n844;
  assign n846 = ~n843 & ~n845;
  assign n847 = ~n841 & n846;
  assign n848 = ~n839 & n847;
  assign n849 = ~n142 & n848;
  assign n850 = n132 & n849;
  assign n851 = ~n837 & n850;
  assign n852 = ~G14gat & ~n851;
  assign n853 = G60gat & G66gat;
  assign n854 = G50gat & n853;
  assign n855 = G56gat & ~n854;
  assign n856 = G47gat & G53gat;
  assign n857 = G37gat & n856;
  assign n858 = G43gat & ~n857;
  assign n859 = G34gat & G40gat;
  assign n860 = G24gat & n859;
  assign n861 = G30gat & ~n860;
  assign n862 = n160 & ~n861;
  assign n863 = ~n858 & n862;
  assign n864 = ~n855 & n863;
  assign n865 = G86gat & G92gat;
  assign n866 = G76gat & n865;
  assign n867 = G82gat & ~n866;
  assign n868 = G73gat & G79gat;
  assign n869 = G63gat & n868;
  assign n870 = G69gat & ~n869;
  assign n871 = ~n867 & ~n870;
  assign n872 = n864 & n871;
  assign n873 = G27gat & n872;
  assign n874 = G14gat & ~n873;
  assign n875 = ~n852 & ~n874;
  assign n876 = G8gat & ~n875;
  assign n877 = ~n835 & ~n876;
  assign n878 = G21gat & n877;
  assign n879 = G27gat & n832;
  assign n880 = G14gat & ~n879;
  assign n881 = ~G8gat & ~n813;
  assign n882 = ~n880 & n881;
  assign n883 = ~G21gat & n882;
  assign n884 = ~n878 & ~n883;
  assign n885 = G11gat & ~n884;
  assign n886 = G17gat & n885;
  assign n887 = G14gat & ~n872;
  assign n888 = ~n852 & ~n887;
  assign n889 = G8gat & ~n888;
  assign n890 = ~n835 & ~n889;
  assign n891 = ~G17gat & n890;
  assign n892 = ~n886 & ~n891;
  assign n893 = G1gat & ~n892;
  assign n894 = ~G8gat & ~n666;
  assign n895 = n174 & ~n865;
  assign n896 = ~G24gat & ~n859;
  assign n897 = G30gat & n896;
  assign n898 = ~n895 & ~n897;
  assign n899 = G99gat & G105gat;
  assign n900 = n173 & ~n899;
  assign n901 = n898 & ~n900;
  assign n902 = ~n77 & n901;
  assign n903 = n172 & ~n856;
  assign n904 = n902 & ~n903;
  assign n905 = ~n434 & n904;
  assign n906 = n178 & ~n853;
  assign n907 = n905 & ~n906;
  assign n908 = n177 & ~n868;
  assign n909 = n907 & ~n908;
  assign n910 = G8gat & ~n909;
  assign n911 = ~n894 & ~n910;
  assign n912 = ~n171 & ~n911;
  assign n913 = G21gat & n894;
  assign n914 = ~n912 & ~n913;
  assign n915 = G27gat & n909;
  assign n916 = G8gat & ~n915;
  assign n917 = ~n668 & ~n916;
  assign n918 = n171 & ~n917;
  assign n919 = n914 & ~n918;
  assign n920 = G14gat & ~n919;
  assign n921 = G95gat & n203;
  assign n922 = ~G34gat & n182;
  assign n923 = ~n921 & ~n922;
  assign n924 = ~n311 & n923;
  assign n925 = ~n295 & n924;
  assign n926 = ~n327 & n925;
  assign n927 = ~n281 & n926;
  assign n928 = ~n73 & n927;
  assign n929 = ~G14gat & ~n928;
  assign n930 = ~n359 & ~n929;
  assign n931 = G8gat & ~n930;
  assign n932 = ~n920 & ~n931;
  assign n933 = ~G1gat & n932;
  assign n934 = ~n893 & ~n933;
  assign n935 = G4gat & n934;
  assign n936 = ~n812 & ~n935;
  assign n937 = keyinput3_G421gat & ~n936;
  assign n938 = ~n804 & ~n937;
  assign n939 = keyinput2_G421gat & ~n938;
  assign n940 = ~n803 & ~n939;
  assign n941 = keyinput1_G421gat & ~n940;
  assign n942 = ~n799 & ~n941;
  assign n943 = keyinput0_G421gat & ~n942;
  assign G421gat = n789 | n943;
  assign n945 = ~keyinput0_G430gat & ~n73;
  assign n946 = keyinput0_G430gat & n104;
  assign n947 = ~n945 & ~n946;
  assign n948 = ~keyinput1_G430gat & ~n947;
  assign n949 = ~G105gat & ~keyinput0_G430gat;
  assign n950 = n74 & ~n949;
  assign n951 = keyinput1_G430gat & ~n950;
  assign n952 = ~n948 & ~n951;
  assign n953 = ~keyinput2_G430gat & ~n952;
  assign n954 = ~keyinput0_G430gat & ~n396;
  assign n955 = keyinput0_G430gat & ~n180;
  assign n956 = ~n954 & ~n955;
  assign n957 = ~keyinput1_G430gat & ~n956;
  assign n958 = keyinput0_G430gat & n72;
  assign n959 = ~keyinput0_G430gat & ~n132;
  assign n960 = ~n958 & ~n959;
  assign n961 = keyinput1_G430gat & ~n960;
  assign n962 = ~n957 & ~n961;
  assign n963 = keyinput2_G430gat & ~n962;
  assign n964 = ~n953 & ~n963;
  assign n965 = ~keyinput3_G430gat & ~n964;
  assign n966 = ~keyinput0_G430gat & n114;
  assign n967 = keyinput0_G430gat & ~n176;
  assign n968 = ~n966 & ~n967;
  assign n969 = ~keyinput1_G430gat & ~n968;
  assign n970 = ~keyinput0_G430gat & n112;
  assign n971 = ~n958 & ~n970;
  assign n972 = keyinput1_G430gat & n971;
  assign n973 = ~n969 & ~n972;
  assign n974 = ~keyinput2_G430gat & ~n973;
  assign n975 = ~keyinput0_G430gat & ~n202;
  assign n976 = ~n958 & ~n975;
  assign n977 = ~keyinput1_G430gat & ~n976;
  assign n978 = ~G108gat & ~keyinput0_G430gat;
  assign n979 = ~n525 & ~n571;
  assign n980 = ~n618 & n979;
  assign n981 = G40gat & n980;
  assign n982 = ~G34gat & ~n981;
  assign n983 = ~n73 & ~n921;
  assign n984 = ~n281 & n983;
  assign n985 = ~n295 & n984;
  assign n986 = ~n311 & ~n985;
  assign n987 = G66gat & ~n525;
  assign n988 = n311 & n987;
  assign n989 = ~n986 & ~n988;
  assign n990 = ~n327 & ~n989;
  assign n991 = G53gat & n979;
  assign n992 = n327 & n991;
  assign n993 = ~n990 & ~n992;
  assign n994 = ~G40gat & n993;
  assign n995 = ~G60gat & ~n987;
  assign n996 = ~G66gat & n985;
  assign n997 = ~n94 & ~n900;
  assign n998 = ~n895 & n997;
  assign n999 = ~n908 & n998;
  assign n1000 = G66gat & n999;
  assign n1001 = ~n996 & ~n1000;
  assign n1002 = G60gat & ~n1001;
  assign n1003 = ~n995 & ~n1002;
  assign n1004 = ~G50gat & ~n1003;
  assign n1005 = G56gat & n1004;
  assign n1006 = ~n178 & n999;
  assign n1007 = ~n1005 & ~n1006;
  assign n1008 = ~n172 & ~n1007;
  assign n1009 = ~G47gat & ~n991;
  assign n1010 = ~G53gat & n989;
  assign n1011 = G53gat & ~n1007;
  assign n1012 = ~n1010 & ~n1011;
  assign n1013 = G47gat & ~n1012;
  assign n1014 = ~n1009 & ~n1013;
  assign n1015 = ~G37gat & ~n1014;
  assign n1016 = G43gat & n1015;
  assign n1017 = ~n1008 & ~n1016;
  assign n1018 = G40gat & ~n1017;
  assign n1019 = ~n994 & ~n1018;
  assign n1020 = G34gat & ~n1019;
  assign n1021 = ~n982 & ~n1020;
  assign n1022 = ~G24gat & ~n1021;
  assign n1023 = ~n837 & ~n839;
  assign n1024 = n143 & n1023;
  assign n1025 = ~G56gat & n1024;
  assign n1026 = n176 & ~n177;
  assign n1027 = ~G66gat & n1026;
  assign n1028 = ~n103 & ~n819;
  assign n1029 = n818 & n1028;
  assign n1030 = G66gat & n1029;
  assign n1031 = ~n1027 & ~n1030;
  assign n1032 = ~G60gat & ~n1031;
  assign n1033 = G60gat & n1024;
  assign n1034 = ~n1032 & ~n1033;
  assign n1035 = G50gat & ~n1034;
  assign n1036 = ~n1004 & ~n1035;
  assign n1037 = G56gat & ~n1036;
  assign n1038 = ~n1025 & ~n1037;
  assign n1039 = ~G43gat & ~n1038;
  assign n1040 = G47gat & ~n1038;
  assign n1041 = ~n178 & n1026;
  assign n1042 = ~n1005 & ~n1041;
  assign n1043 = ~G53gat & n1042;
  assign n1044 = ~G47gat & ~n1043;
  assign n1045 = ~G56gat & n1029;
  assign n1046 = G60gat & n1029;
  assign n1047 = ~n1032 & ~n1046;
  assign n1048 = G50gat & ~n1047;
  assign n1049 = ~n1004 & ~n1048;
  assign n1050 = G56gat & ~n1049;
  assign n1051 = ~n1045 & ~n1050;
  assign n1052 = G53gat & n1051;
  assign n1053 = n1044 & ~n1052;
  assign n1054 = ~n1040 & ~n1053;
  assign n1055 = G37gat & ~n1054;
  assign n1056 = ~n1015 & ~n1055;
  assign n1057 = G43gat & ~n1056;
  assign n1058 = ~n1039 & ~n1057;
  assign n1059 = ~G40gat & ~n1058;
  assign n1060 = n160 & n871;
  assign n1061 = ~G56gat & n1060;
  assign n1062 = ~G66gat & n1024;
  assign n1063 = G66gat & n1060;
  assign n1064 = ~n1062 & ~n1063;
  assign n1065 = G60gat & ~n1064;
  assign n1066 = ~n1032 & ~n1065;
  assign n1067 = G50gat & ~n1066;
  assign n1068 = ~n1004 & ~n1067;
  assign n1069 = G56gat & ~n1068;
  assign n1070 = ~n1061 & ~n1069;
  assign n1071 = ~G43gat & ~n1070;
  assign n1072 = ~G53gat & ~n1038;
  assign n1073 = G53gat & ~n1070;
  assign n1074 = ~n1072 & ~n1073;
  assign n1075 = G47gat & ~n1074;
  assign n1076 = ~n1053 & ~n1075;
  assign n1077 = G37gat & ~n1076;
  assign n1078 = ~n1015 & ~n1077;
  assign n1079 = G43gat & ~n1078;
  assign n1080 = ~n1071 & ~n1079;
  assign n1081 = G40gat & ~n1080;
  assign n1082 = ~n1059 & ~n1081;
  assign n1083 = G34gat & ~n1082;
  assign n1084 = ~n172 & ~n1042;
  assign n1085 = ~n1016 & ~n1084;
  assign n1086 = ~G40gat & n1085;
  assign n1087 = ~G34gat & ~n1086;
  assign n1088 = ~G43gat & ~n1051;
  assign n1089 = G47gat & ~n1051;
  assign n1090 = ~n1053 & ~n1089;
  assign n1091 = G37gat & ~n1090;
  assign n1092 = ~n1015 & ~n1091;
  assign n1093 = G43gat & ~n1092;
  assign n1094 = ~n1088 & ~n1093;
  assign n1095 = G40gat & n1094;
  assign n1096 = n1087 & ~n1095;
  assign n1097 = ~n1083 & ~n1096;
  assign n1098 = G24gat & ~n1097;
  assign n1099 = ~n1022 & ~n1098;
  assign n1100 = G30gat & ~n1099;
  assign n1101 = ~G43gat & n1069;
  assign n1102 = ~n1079 & ~n1101;
  assign n1103 = ~G30gat & ~n1102;
  assign n1104 = ~n1100 & ~n1103;
  assign n1105 = ~G17gat & ~n1104;
  assign n1106 = G30gat & n1022;
  assign n1107 = ~n182 & ~n1085;
  assign n1108 = ~n1106 & ~n1107;
  assign n1109 = ~G27gat & ~n1108;
  assign n1110 = ~G30gat & ~n1094;
  assign n1111 = G34gat & ~n1094;
  assign n1112 = ~n1096 & ~n1111;
  assign n1113 = G24gat & ~n1112;
  assign n1114 = ~n1022 & ~n1113;
  assign n1115 = G30gat & ~n1114;
  assign n1116 = ~n1110 & ~n1115;
  assign n1117 = G27gat & ~n1116;
  assign n1118 = ~n1109 & ~n1117;
  assign n1119 = ~G21gat & ~n1118;
  assign n1120 = ~G30gat & ~n1058;
  assign n1121 = G34gat & ~n1058;
  assign n1122 = ~n1096 & ~n1121;
  assign n1123 = G24gat & ~n1122;
  assign n1124 = ~n1022 & ~n1123;
  assign n1125 = G30gat & ~n1124;
  assign n1126 = ~n1120 & ~n1125;
  assign n1127 = ~G27gat & ~n1126;
  assign n1128 = ~G30gat & ~n1080;
  assign n1129 = ~n1100 & ~n1128;
  assign n1130 = G27gat & ~n1129;
  assign n1131 = ~n1127 & ~n1130;
  assign n1132 = G21gat & ~n1131;
  assign n1133 = ~n1119 & ~n1132;
  assign n1134 = G11gat & ~n1133;
  assign n1135 = G27gat & n980;
  assign n1136 = ~n665 & n1135;
  assign n1137 = ~G21gat & n1136;
  assign n1138 = ~G11gat & ~n1137;
  assign n1139 = ~n343 & ~n993;
  assign n1140 = n343 & n981;
  assign n1141 = ~n1139 & ~n1140;
  assign n1142 = ~G27gat & n1141;
  assign n1143 = ~n182 & ~n1017;
  assign n1144 = ~n1106 & ~n1143;
  assign n1145 = G27gat & ~n1144;
  assign n1146 = ~n1142 & ~n1145;
  assign n1147 = G21gat & n1146;
  assign n1148 = n1138 & ~n1147;
  assign n1149 = ~n1134 & ~n1148;
  assign n1150 = G17gat & ~n1149;
  assign n1151 = ~n1105 & ~n1150;
  assign n1152 = ~G4gat & ~n1151;
  assign n1153 = ~n571 & ~n665;
  assign n1154 = ~n618 & n1153;
  assign n1155 = ~G14gat & ~n1154;
  assign n1156 = n172 & n1009;
  assign n1157 = ~G47gat & n172;
  assign n1158 = n995 & ~n1157;
  assign n1159 = n178 & n1158;
  assign n1160 = ~n1156 & ~n1159;
  assign n1161 = ~n922 & n1160;
  assign n1162 = G14gat & ~n1161;
  assign n1163 = ~n1140 & n1162;
  assign n1164 = ~n1155 & ~n1163;
  assign n1165 = ~G8gat & n1164;
  assign n1166 = G60gat & n996;
  assign n1167 = ~n995 & ~n1166;
  assign n1168 = n178 & ~n1167;
  assign n1169 = ~n172 & n1168;
  assign n1170 = G53gat & n1168;
  assign n1171 = ~n1010 & ~n1170;
  assign n1172 = G47gat & ~n1171;
  assign n1173 = ~n1009 & ~n1172;
  assign n1174 = n172 & ~n1173;
  assign n1175 = ~n1169 & ~n1174;
  assign n1176 = ~n182 & n1175;
  assign n1177 = G40gat & ~n1175;
  assign n1178 = ~n994 & ~n1177;
  assign n1179 = G34gat & ~n1178;
  assign n1180 = ~n982 & ~n1179;
  assign n1181 = n182 & n1180;
  assign n1182 = ~n1176 & ~n1181;
  assign n1183 = ~G14gat & n1182;
  assign n1184 = ~n172 & n1005;
  assign n1185 = ~n1016 & ~n1184;
  assign n1186 = ~n182 & ~n1185;
  assign n1187 = ~n1106 & ~n1186;
  assign n1188 = G14gat & ~n1187;
  assign n1189 = ~n1183 & ~n1188;
  assign n1190 = G8gat & n1189;
  assign n1191 = ~n1165 & ~n1190;
  assign n1192 = ~n171 & ~n1191;
  assign n1193 = G27gat & n1182;
  assign n1194 = ~n1142 & ~n1193;
  assign n1195 = ~G14gat & ~n1194;
  assign n1196 = G14gat & ~n1146;
  assign n1197 = ~n1195 & ~n1196;
  assign n1198 = G21gat & n1197;
  assign n1199 = ~n1137 & ~n1198;
  assign n1200 = G8gat & ~n1199;
  assign n1201 = G27gat & n1154;
  assign n1202 = ~G14gat & ~n1201;
  assign n1203 = G14gat & ~n1136;
  assign n1204 = ~n1202 & ~n1203;
  assign n1205 = ~G21gat & ~n1204;
  assign n1206 = G21gat & ~n1164;
  assign n1207 = ~n1205 & ~n1206;
  assign n1208 = ~G8gat & n1207;
  assign n1209 = ~n1200 & ~n1208;
  assign n1210 = n171 & ~n1209;
  assign n1211 = ~n1192 & ~n1210;
  assign n1212 = ~G1gat & n1211;
  assign n1213 = G50gat & ~G60gat;
  assign n1214 = n1027 & n1213;
  assign n1215 = ~n1004 & ~n1214;
  assign n1216 = G56gat & ~n1215;
  assign n1217 = ~G43gat & n1216;
  assign n1218 = ~n617 & ~n1216;
  assign n1219 = ~G47gat & n1043;
  assign n1220 = ~n1218 & ~n1219;
  assign n1221 = G37gat & n1220;
  assign n1222 = ~n1015 & ~n1221;
  assign n1223 = G43gat & ~n1222;
  assign n1224 = ~n1217 & ~n1223;
  assign n1225 = ~G30gat & ~n1224;
  assign n1226 = ~n664 & n1224;
  assign n1227 = ~G34gat & n1086;
  assign n1228 = ~n1226 & ~n1227;
  assign n1229 = G24gat & n1228;
  assign n1230 = ~n1022 & ~n1229;
  assign n1231 = G30gat & ~n1230;
  assign n1232 = ~n1225 & ~n1231;
  assign n1233 = ~G14gat & ~n1232;
  assign n1234 = G50gat & n1032;
  assign n1235 = ~n1004 & ~n1234;
  assign n1236 = G56gat & ~n1235;
  assign n1237 = ~G43gat & n1236;
  assign n1238 = G47gat & n1236;
  assign n1239 = ~n1053 & ~n1238;
  assign n1240 = G37gat & ~n1239;
  assign n1241 = ~n1015 & ~n1240;
  assign n1242 = G43gat & ~n1241;
  assign n1243 = ~n1237 & ~n1242;
  assign n1244 = ~G30gat & ~n1243;
  assign n1245 = G34gat & ~n1243;
  assign n1246 = ~n1096 & ~n1245;
  assign n1247 = G24gat & ~n1246;
  assign n1248 = ~n1022 & ~n1247;
  assign n1249 = G30gat & ~n1248;
  assign n1250 = ~n1244 & ~n1249;
  assign n1251 = G14gat & ~n1250;
  assign n1252 = ~n1233 & ~n1251;
  assign n1253 = ~G8gat & ~n1252;
  assign n1254 = G60gat & n1062;
  assign n1255 = ~n1032 & ~n1254;
  assign n1256 = G50gat & ~n1255;
  assign n1257 = ~n1004 & ~n1256;
  assign n1258 = G56gat & ~n1257;
  assign n1259 = ~G43gat & n1258;
  assign n1260 = G53gat & n1258;
  assign n1261 = ~n1072 & ~n1260;
  assign n1262 = G47gat & ~n1261;
  assign n1263 = ~n1053 & ~n1262;
  assign n1264 = G37gat & ~n1263;
  assign n1265 = ~n1015 & ~n1264;
  assign n1266 = G43gat & ~n1265;
  assign n1267 = ~n1259 & ~n1266;
  assign n1268 = ~G30gat & ~n1267;
  assign n1269 = G40gat & ~n1267;
  assign n1270 = ~n1059 & ~n1269;
  assign n1271 = G34gat & ~n1270;
  assign n1272 = ~n1096 & ~n1271;
  assign n1273 = G24gat & ~n1272;
  assign n1274 = ~n1022 & ~n1273;
  assign n1275 = G30gat & ~n1274;
  assign n1276 = ~n1268 & ~n1275;
  assign n1277 = ~G14gat & ~n1276;
  assign n1278 = G14gat & ~n1104;
  assign n1279 = ~n1277 & ~n1278;
  assign n1280 = G8gat & ~n1279;
  assign n1281 = ~n1253 & ~n1280;
  assign n1282 = ~G17gat & ~n1281;
  assign n1283 = G21gat & ~n1252;
  assign n1284 = G14gat & ~n1116;
  assign n1285 = ~n1233 & ~n1284;
  assign n1286 = G27gat & ~n1285;
  assign n1287 = ~n1109 & ~n1286;
  assign n1288 = ~G21gat & ~n1287;
  assign n1289 = ~n1283 & ~n1288;
  assign n1290 = ~G8gat & ~n1289;
  assign n1291 = G14gat & ~n1129;
  assign n1292 = ~n1277 & ~n1291;
  assign n1293 = G27gat & ~n1292;
  assign n1294 = ~n1127 & ~n1293;
  assign n1295 = G21gat & ~n1294;
  assign n1296 = ~n1119 & ~n1295;
  assign n1297 = G8gat & ~n1296;
  assign n1298 = ~n1290 & ~n1297;
  assign n1299 = G11gat & ~n1298;
  assign n1300 = ~n1148 & ~n1299;
  assign n1301 = G17gat & ~n1300;
  assign n1302 = ~n1282 & ~n1301;
  assign n1303 = G1gat & ~n1302;
  assign n1304 = ~n1212 & ~n1303;
  assign n1305 = G4gat & ~n1304;
  assign n1306 = ~n1152 & ~n1305;
  assign n1307 = keyinput0_G430gat & ~n1306;
  assign n1308 = ~n978 & ~n1307;
  assign n1309 = keyinput1_G430gat & ~n1308;
  assign n1310 = ~n977 & ~n1309;
  assign n1311 = keyinput2_G430gat & ~n1310;
  assign n1312 = ~n974 & ~n1311;
  assign n1313 = keyinput3_G430gat & ~n1312;
  assign G430gat = n965 | n1313;
  assign n1315 = ~keyinput0_G431gat & ~n73;
  assign n1316 = keyinput0_G431gat & n104;
  assign n1317 = ~n1315 & ~n1316;
  assign n1318 = ~keyinput1_G431gat & ~n1317;
  assign n1319 = ~G105gat & ~keyinput0_G431gat;
  assign n1320 = n74 & ~n1319;
  assign n1321 = keyinput1_G431gat & ~n1320;
  assign n1322 = ~n1318 & ~n1321;
  assign n1323 = ~keyinput2_G431gat & ~n1322;
  assign n1324 = ~keyinput0_G431gat & ~n396;
  assign n1325 = keyinput0_G431gat & ~n180;
  assign n1326 = ~n1324 & ~n1325;
  assign n1327 = ~keyinput1_G431gat & ~n1326;
  assign n1328 = keyinput0_G431gat & n72;
  assign n1329 = ~keyinput0_G431gat & ~n132;
  assign n1330 = ~n1328 & ~n1329;
  assign n1331 = keyinput1_G431gat & ~n1330;
  assign n1332 = ~n1327 & ~n1331;
  assign n1333 = keyinput2_G431gat & ~n1332;
  assign n1334 = ~n1323 & ~n1333;
  assign n1335 = ~keyinput3_G431gat & ~n1334;
  assign n1336 = ~keyinput0_G431gat & n114;
  assign n1337 = keyinput0_G431gat & ~n176;
  assign n1338 = ~n1336 & ~n1337;
  assign n1339 = ~keyinput1_G431gat & ~n1338;
  assign n1340 = ~keyinput0_G431gat & n112;
  assign n1341 = ~n1328 & ~n1340;
  assign n1342 = keyinput1_G431gat & n1341;
  assign n1343 = ~n1339 & ~n1342;
  assign n1344 = ~keyinput2_G431gat & ~n1343;
  assign n1345 = ~keyinput0_G431gat & ~n202;
  assign n1346 = ~n1328 & ~n1345;
  assign n1347 = ~keyinput1_G431gat & ~n1346;
  assign n1348 = ~G108gat & ~keyinput0_G431gat;
  assign n1349 = ~n431 & ~n477;
  assign n1350 = ~n524 & n1349;
  assign n1351 = ~n571 & ~n1350;
  assign n1352 = ~n618 & n1351;
  assign n1353 = G40gat & ~n1352;
  assign n1354 = ~G34gat & ~n1353;
  assign n1355 = ~G73gat & n177;
  assign n1356 = G92gat & ~n431;
  assign n1357 = n281 & ~n1356;
  assign n1358 = ~n984 & ~n1357;
  assign n1359 = ~n1355 & ~n1358;
  assign n1360 = G79gat & n1349;
  assign n1361 = n295 & ~n1360;
  assign n1362 = ~n1359 & ~n1361;
  assign n1363 = ~n311 & ~n1362;
  assign n1364 = ~n477 & ~n524;
  assign n1365 = G66gat & ~n1364;
  assign n1366 = n311 & n1365;
  assign n1367 = ~n1363 & ~n1366;
  assign n1368 = ~n327 & ~n1367;
  assign n1369 = ~n571 & ~n1364;
  assign n1370 = G53gat & n1369;
  assign n1371 = n327 & n1370;
  assign n1372 = ~n1368 & ~n1371;
  assign n1373 = ~G40gat & ~n1372;
  assign n1374 = ~G86gat & ~n1356;
  assign n1375 = G92gat & n997;
  assign n1376 = ~G92gat & n983;
  assign n1377 = ~n1375 & ~n1376;
  assign n1378 = G86gat & ~n1377;
  assign n1379 = ~n1374 & ~n1378;
  assign n1380 = ~G76gat & ~n1379;
  assign n1381 = G82gat & n1380;
  assign n1382 = ~n174 & n997;
  assign n1383 = ~n1381 & ~n1382;
  assign n1384 = ~n908 & n1383;
  assign n1385 = ~n906 & ~n1384;
  assign n1386 = ~G73gat & ~n1360;
  assign n1387 = ~G79gat & ~n1358;
  assign n1388 = ~n868 & ~n1387;
  assign n1389 = ~n1386 & n1388;
  assign n1390 = n177 & n1389;
  assign n1391 = n1385 & ~n1390;
  assign n1392 = ~G60gat & n1365;
  assign n1393 = ~n295 & n1374;
  assign n1394 = n174 & n1393;
  assign n1395 = ~n1361 & ~n1394;
  assign n1396 = ~G66gat & ~n1395;
  assign n1397 = G60gat & n1396;
  assign n1398 = ~n1392 & ~n1397;
  assign n1399 = n178 & ~n1398;
  assign n1400 = ~n1391 & ~n1399;
  assign n1401 = ~n903 & ~n1400;
  assign n1402 = ~G47gat & n1370;
  assign n1403 = ~n311 & ~n1395;
  assign n1404 = ~n1366 & ~n1403;
  assign n1405 = ~G53gat & ~n1404;
  assign n1406 = G47gat & n1405;
  assign n1407 = ~n1402 & ~n1406;
  assign n1408 = n172 & ~n1407;
  assign n1409 = ~n1401 & ~n1408;
  assign n1410 = G40gat & ~n1409;
  assign n1411 = ~n1373 & ~n1410;
  assign n1412 = G34gat & ~n1411;
  assign n1413 = ~n1354 & ~n1412;
  assign n1414 = ~G24gat & ~n1413;
  assign n1415 = ~n1374 & ~n1376;
  assign n1416 = n174 & ~n1415;
  assign n1417 = ~n908 & ~n1416;
  assign n1418 = ~n1390 & ~n1417;
  assign n1419 = G66gat & n1418;
  assign n1420 = ~n1396 & ~n1419;
  assign n1421 = G60gat & ~n1420;
  assign n1422 = ~n1392 & ~n1421;
  assign n1423 = ~G50gat & ~n1422;
  assign n1424 = G56gat & n1423;
  assign n1425 = ~n178 & n1418;
  assign n1426 = ~n1424 & ~n1425;
  assign n1427 = G53gat & ~n1426;
  assign n1428 = ~n1405 & ~n1427;
  assign n1429 = G47gat & ~n1428;
  assign n1430 = ~n1402 & ~n1429;
  assign n1431 = ~G37gat & ~n1430;
  assign n1432 = G43gat & n1431;
  assign n1433 = ~n174 & n270;
  assign n1434 = ~n1381 & ~n1433;
  assign n1435 = ~n177 & ~n1434;
  assign n1436 = G79gat & ~n1383;
  assign n1437 = ~n1387 & ~n1436;
  assign n1438 = G73gat & ~n1437;
  assign n1439 = ~n1386 & ~n1438;
  assign n1440 = ~G63gat & ~n1439;
  assign n1441 = G69gat & n1440;
  assign n1442 = ~n1435 & ~n1441;
  assign n1443 = ~n178 & ~n1442;
  assign n1444 = ~n1424 & ~n1443;
  assign n1445 = ~n172 & ~n1444;
  assign n1446 = ~n1432 & ~n1445;
  assign n1447 = ~G40gat & ~n1446;
  assign n1448 = ~G82gat & n1028;
  assign n1449 = G86gat & n1028;
  assign n1450 = G92gat & n1028;
  assign n1451 = ~G92gat & n270;
  assign n1452 = ~n1450 & ~n1451;
  assign n1453 = ~G86gat & ~n1452;
  assign n1454 = ~n1449 & ~n1453;
  assign n1455 = G76gat & ~n1454;
  assign n1456 = ~n1380 & ~n1455;
  assign n1457 = G82gat & ~n1456;
  assign n1458 = ~n1448 & ~n1457;
  assign n1459 = ~G69gat & ~n1458;
  assign n1460 = G73gat & ~n1458;
  assign n1461 = ~G79gat & n1434;
  assign n1462 = ~G73gat & ~n1461;
  assign n1463 = G79gat & n1458;
  assign n1464 = n1462 & ~n1463;
  assign n1465 = ~n1460 & ~n1464;
  assign n1466 = G63gat & ~n1465;
  assign n1467 = ~n1440 & ~n1466;
  assign n1468 = G69gat & ~n1467;
  assign n1469 = ~n1459 & ~n1468;
  assign n1470 = ~G56gat & ~n1469;
  assign n1471 = ~n820 & ~n1469;
  assign n1472 = ~n177 & n1381;
  assign n1473 = ~n1441 & ~n1472;
  assign n1474 = ~G66gat & ~n1473;
  assign n1475 = ~G60gat & n1474;
  assign n1476 = ~n1471 & ~n1475;
  assign n1477 = G50gat & ~n1476;
  assign n1478 = ~n1423 & ~n1477;
  assign n1479 = G56gat & ~n1478;
  assign n1480 = ~n1470 & ~n1479;
  assign n1481 = ~G43gat & ~n1480;
  assign n1482 = ~n617 & n1480;
  assign n1483 = ~n178 & ~n1473;
  assign n1484 = ~n1424 & ~n1483;
  assign n1485 = n617 & n1484;
  assign n1486 = ~n1482 & ~n1485;
  assign n1487 = G37gat & n1486;
  assign n1488 = ~n1431 & ~n1487;
  assign n1489 = G43gat & ~n1488;
  assign n1490 = ~n1481 & ~n1489;
  assign n1491 = G40gat & ~n1490;
  assign n1492 = ~n1447 & ~n1491;
  assign n1493 = ~G34gat & ~n1492;
  assign n1494 = ~G82gat & n143;
  assign n1495 = G86gat & n143;
  assign n1496 = ~n1453 & ~n1495;
  assign n1497 = G76gat & ~n1496;
  assign n1498 = ~n1380 & ~n1497;
  assign n1499 = G82gat & ~n1498;
  assign n1500 = ~n1494 & ~n1499;
  assign n1501 = ~G69gat & ~n1500;
  assign n1502 = G73gat & ~n1500;
  assign n1503 = ~n1464 & ~n1502;
  assign n1504 = G63gat & ~n1503;
  assign n1505 = ~n1440 & ~n1504;
  assign n1506 = G69gat & ~n1505;
  assign n1507 = ~n1501 & ~n1506;
  assign n1508 = ~G56gat & ~n1507;
  assign n1509 = G76gat & ~G86gat;
  assign n1510 = n1451 & n1509;
  assign n1511 = ~n1380 & ~n1510;
  assign n1512 = G82gat & ~n1511;
  assign n1513 = ~G69gat & n1512;
  assign n1514 = ~n523 & ~n1512;
  assign n1515 = ~G73gat & n1461;
  assign n1516 = ~n1514 & ~n1515;
  assign n1517 = G63gat & n1516;
  assign n1518 = ~n1440 & ~n1517;
  assign n1519 = G69gat & ~n1518;
  assign n1520 = ~n1513 & ~n1519;
  assign n1521 = G66gat & ~n1520;
  assign n1522 = ~n1474 & ~n1521;
  assign n1523 = ~G60gat & ~n1522;
  assign n1524 = G60gat & ~n1507;
  assign n1525 = ~n1523 & ~n1524;
  assign n1526 = G50gat & ~n1525;
  assign n1527 = ~n1423 & ~n1526;
  assign n1528 = G56gat & ~n1527;
  assign n1529 = ~n1508 & ~n1528;
  assign n1530 = ~G43gat & ~n1529;
  assign n1531 = ~G53gat & ~n1484;
  assign n1532 = n1213 & n1474;
  assign n1533 = ~n1423 & ~n1532;
  assign n1534 = G56gat & ~n1533;
  assign n1535 = ~n822 & ~n1520;
  assign n1536 = ~n1534 & ~n1535;
  assign n1537 = G53gat & ~n1536;
  assign n1538 = ~n1531 & ~n1537;
  assign n1539 = ~G47gat & ~n1538;
  assign n1540 = G47gat & ~n1529;
  assign n1541 = ~n1539 & ~n1540;
  assign n1542 = G37gat & ~n1541;
  assign n1543 = ~n1431 & ~n1542;
  assign n1544 = G43gat & ~n1543;
  assign n1545 = ~n1530 & ~n1544;
  assign n1546 = ~G40gat & ~n1545;
  assign n1547 = ~G82gat & n160;
  assign n1548 = G92gat & n160;
  assign n1549 = ~G92gat & n143;
  assign n1550 = ~n1548 & ~n1549;
  assign n1551 = G86gat & ~n1550;
  assign n1552 = ~n1453 & ~n1551;
  assign n1553 = G76gat & ~n1552;
  assign n1554 = ~n1380 & ~n1553;
  assign n1555 = G82gat & ~n1554;
  assign n1556 = ~n1547 & ~n1555;
  assign n1557 = ~G69gat & ~n1556;
  assign n1558 = ~G79gat & ~n1500;
  assign n1559 = G79gat & ~n1556;
  assign n1560 = ~n1558 & ~n1559;
  assign n1561 = G73gat & ~n1560;
  assign n1562 = ~n1464 & ~n1561;
  assign n1563 = G63gat & ~n1562;
  assign n1564 = ~n1440 & ~n1563;
  assign n1565 = G69gat & ~n1564;
  assign n1566 = ~n1557 & ~n1565;
  assign n1567 = ~G56gat & ~n1566;
  assign n1568 = G76gat & n1453;
  assign n1569 = ~n1380 & ~n1568;
  assign n1570 = G82gat & ~n1569;
  assign n1571 = ~G69gat & n1570;
  assign n1572 = G73gat & n1570;
  assign n1573 = ~n1464 & ~n1572;
  assign n1574 = G63gat & ~n1573;
  assign n1575 = ~n1440 & ~n1574;
  assign n1576 = G69gat & ~n1575;
  assign n1577 = ~n1571 & ~n1576;
  assign n1578 = ~G66gat & ~n1577;
  assign n1579 = G66gat & ~n1566;
  assign n1580 = ~n1578 & ~n1579;
  assign n1581 = G60gat & ~n1580;
  assign n1582 = ~n1523 & ~n1581;
  assign n1583 = G50gat & ~n1582;
  assign n1584 = ~n1423 & ~n1583;
  assign n1585 = G56gat & ~n1584;
  assign n1586 = ~n1567 & ~n1585;
  assign n1587 = ~G43gat & ~n1586;
  assign n1588 = ~G56gat & ~n1577;
  assign n1589 = G60gat & ~n1577;
  assign n1590 = ~n1523 & ~n1589;
  assign n1591 = G50gat & ~n1590;
  assign n1592 = ~n1423 & ~n1591;
  assign n1593 = G56gat & ~n1592;
  assign n1594 = ~n1588 & ~n1593;
  assign n1595 = ~G53gat & ~n1594;
  assign n1596 = G53gat & ~n1586;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = G47gat & ~n1597;
  assign n1599 = ~n1539 & ~n1598;
  assign n1600 = G37gat & ~n1599;
  assign n1601 = ~n1431 & ~n1600;
  assign n1602 = G43gat & ~n1601;
  assign n1603 = ~n1587 & ~n1602;
  assign n1604 = G40gat & ~n1603;
  assign n1605 = ~n1546 & ~n1604;
  assign n1606 = G34gat & ~n1605;
  assign n1607 = ~n1493 & ~n1606;
  assign n1608 = G24gat & ~n1607;
  assign n1609 = ~n1414 & ~n1608;
  assign n1610 = G30gat & ~n1609;
  assign n1611 = G86gat & n1549;
  assign n1612 = ~n1453 & ~n1611;
  assign n1613 = G76gat & ~n1612;
  assign n1614 = ~n1380 & ~n1613;
  assign n1615 = G82gat & ~n1614;
  assign n1616 = ~G69gat & n1615;
  assign n1617 = G79gat & n1615;
  assign n1618 = ~n1558 & ~n1617;
  assign n1619 = G73gat & ~n1618;
  assign n1620 = ~n1464 & ~n1619;
  assign n1621 = G63gat & ~n1620;
  assign n1622 = ~n1440 & ~n1621;
  assign n1623 = G69gat & ~n1622;
  assign n1624 = ~n1616 & ~n1623;
  assign n1625 = ~G56gat & ~n1624;
  assign n1626 = G66gat & ~n1624;
  assign n1627 = ~n1578 & ~n1626;
  assign n1628 = G60gat & ~n1627;
  assign n1629 = ~n1523 & ~n1628;
  assign n1630 = G50gat & ~n1629;
  assign n1631 = ~n1423 & ~n1630;
  assign n1632 = G56gat & ~n1631;
  assign n1633 = ~n1625 & ~n1632;
  assign n1634 = G53gat & ~n1633;
  assign n1635 = ~n1595 & ~n1634;
  assign n1636 = G47gat & ~n1635;
  assign n1637 = ~n1539 & ~n1636;
  assign n1638 = G37gat & ~n1637;
  assign n1639 = ~n1431 & ~n1638;
  assign n1640 = G43gat & ~n1639;
  assign n1641 = ~G69gat & n1555;
  assign n1642 = ~n1565 & ~n1641;
  assign n1643 = ~G56gat & ~n1642;
  assign n1644 = ~n1632 & ~n1643;
  assign n1645 = ~G43gat & ~n1644;
  assign n1646 = ~n1640 & ~n1645;
  assign n1647 = ~G30gat & ~n1646;
  assign n1648 = ~n1610 & ~n1647;
  assign n1649 = ~G17gat & ~n1648;
  assign n1650 = G27gat & ~n1352;
  assign n1651 = ~n665 & n1650;
  assign n1652 = ~G21gat & ~n1651;
  assign n1653 = ~n343 & n1372;
  assign n1654 = n343 & n1353;
  assign n1655 = ~n1653 & ~n1654;
  assign n1656 = ~G27gat & n1655;
  assign n1657 = G30gat & n1414;
  assign n1658 = ~n182 & ~n1409;
  assign n1659 = ~n1657 & ~n1658;
  assign n1660 = G27gat & ~n1659;
  assign n1661 = ~n1656 & ~n1660;
  assign n1662 = G21gat & ~n1661;
  assign n1663 = ~n1652 & ~n1662;
  assign n1664 = ~G11gat & ~n1663;
  assign n1665 = ~n182 & ~n1446;
  assign n1666 = ~n1657 & ~n1665;
  assign n1667 = ~G27gat & ~n1666;
  assign n1668 = ~G30gat & ~n1490;
  assign n1669 = G34gat & ~n1490;
  assign n1670 = ~n1493 & ~n1669;
  assign n1671 = G24gat & ~n1670;
  assign n1672 = ~n1414 & ~n1671;
  assign n1673 = G30gat & ~n1672;
  assign n1674 = ~n1668 & ~n1673;
  assign n1675 = G27gat & ~n1674;
  assign n1676 = ~n1667 & ~n1675;
  assign n1677 = ~G21gat & ~n1676;
  assign n1678 = ~G30gat & ~n1545;
  assign n1679 = G34gat & ~n1545;
  assign n1680 = ~n1493 & ~n1679;
  assign n1681 = G24gat & ~n1680;
  assign n1682 = ~n1414 & ~n1681;
  assign n1683 = G30gat & ~n1682;
  assign n1684 = ~n1678 & ~n1683;
  assign n1685 = ~G27gat & ~n1684;
  assign n1686 = ~G30gat & ~n1603;
  assign n1687 = ~n1610 & ~n1686;
  assign n1688 = G27gat & ~n1687;
  assign n1689 = ~n1685 & ~n1688;
  assign n1690 = G21gat & ~n1689;
  assign n1691 = ~n1677 & ~n1690;
  assign n1692 = G11gat & ~n1691;
  assign n1693 = ~n1664 & ~n1692;
  assign n1694 = G17gat & ~n1693;
  assign n1695 = ~n1649 & ~n1694;
  assign n1696 = ~G4gat & ~n1695;
  assign n1697 = G24gat & ~G34gat;
  assign n1698 = n1447 & n1697;
  assign n1699 = ~n1414 & ~n1698;
  assign n1700 = G30gat & ~n1699;
  assign n1701 = G37gat & ~G47gat;
  assign n1702 = n1531 & n1701;
  assign n1703 = ~n1431 & ~n1702;
  assign n1704 = G43gat & ~n1703;
  assign n1705 = ~n824 & ~n1536;
  assign n1706 = ~n1704 & ~n1705;
  assign n1707 = ~n826 & ~n1706;
  assign n1708 = ~n1700 & ~n1707;
  assign n1709 = ~G14gat & ~n1708;
  assign n1710 = ~G43gat & ~n1594;
  assign n1711 = G47gat & ~n1594;
  assign n1712 = ~n1539 & ~n1711;
  assign n1713 = G37gat & ~n1712;
  assign n1714 = ~n1431 & ~n1713;
  assign n1715 = G43gat & ~n1714;
  assign n1716 = ~n1710 & ~n1715;
  assign n1717 = ~G30gat & ~n1716;
  assign n1718 = G34gat & ~n1716;
  assign n1719 = ~n1493 & ~n1718;
  assign n1720 = G24gat & ~n1719;
  assign n1721 = ~n1414 & ~n1720;
  assign n1722 = G30gat & ~n1721;
  assign n1723 = ~n1717 & ~n1722;
  assign n1724 = G14gat & ~n1723;
  assign n1725 = ~n1709 & ~n1724;
  assign n1726 = ~G8gat & ~n1725;
  assign n1727 = ~G43gat & ~n1633;
  assign n1728 = ~n1640 & ~n1727;
  assign n1729 = ~G30gat & ~n1728;
  assign n1730 = G40gat & ~n1728;
  assign n1731 = ~n1546 & ~n1730;
  assign n1732 = G34gat & ~n1731;
  assign n1733 = ~n1493 & ~n1732;
  assign n1734 = G24gat & ~n1733;
  assign n1735 = ~n1414 & ~n1734;
  assign n1736 = G30gat & ~n1735;
  assign n1737 = ~n1729 & ~n1736;
  assign n1738 = ~G14gat & ~n1737;
  assign n1739 = G14gat & ~n1648;
  assign n1740 = ~n1738 & ~n1739;
  assign n1741 = G8gat & ~n1740;
  assign n1742 = ~n1726 & ~n1741;
  assign n1743 = ~G17gat & ~n1742;
  assign n1744 = G21gat & ~n1725;
  assign n1745 = G14gat & ~n1674;
  assign n1746 = ~n1709 & ~n1745;
  assign n1747 = G27gat & ~n1746;
  assign n1748 = ~n1667 & ~n1747;
  assign n1749 = ~G21gat & ~n1748;
  assign n1750 = ~n1744 & ~n1749;
  assign n1751 = ~G8gat & ~n1750;
  assign n1752 = G14gat & ~n1687;
  assign n1753 = ~n1738 & ~n1752;
  assign n1754 = G27gat & ~n1753;
  assign n1755 = ~n1685 & ~n1754;
  assign n1756 = G21gat & ~n1755;
  assign n1757 = ~n1677 & ~n1756;
  assign n1758 = G8gat & ~n1757;
  assign n1759 = ~n1751 & ~n1758;
  assign n1760 = G11gat & ~n1759;
  assign n1761 = ~n1664 & ~n1760;
  assign n1762 = G17gat & ~n1761;
  assign n1763 = ~n1743 & ~n1762;
  assign n1764 = G1gat & ~n1763;
  assign n1765 = ~n618 & n1369;
  assign n1766 = ~n665 & ~n1765;
  assign n1767 = ~G14gat & ~n1766;
  assign n1768 = ~n327 & ~n1404;
  assign n1769 = ~n1371 & ~n1768;
  assign n1770 = ~n922 & ~n1769;
  assign n1771 = n182 & n1354;
  assign n1772 = ~n1770 & ~n1771;
  assign n1773 = G14gat & ~n1772;
  assign n1774 = ~n1767 & ~n1773;
  assign n1775 = ~G8gat & ~n1774;
  assign n1776 = ~n903 & ~n1426;
  assign n1777 = ~n1408 & ~n1776;
  assign n1778 = ~n182 & n1777;
  assign n1779 = G40gat & ~n1777;
  assign n1780 = ~n1373 & ~n1779;
  assign n1781 = G34gat & ~n1780;
  assign n1782 = ~n1354 & ~n1781;
  assign n1783 = n182 & n1782;
  assign n1784 = ~n1778 & ~n1783;
  assign n1785 = ~G14gat & n1784;
  assign n1786 = ~n172 & ~n1484;
  assign n1787 = ~n1432 & ~n1786;
  assign n1788 = ~n182 & ~n1787;
  assign n1789 = ~n1657 & ~n1788;
  assign n1790 = G14gat & ~n1789;
  assign n1791 = ~n1785 & ~n1790;
  assign n1792 = G8gat & ~n1791;
  assign n1793 = ~n1775 & ~n1792;
  assign n1794 = ~n171 & ~n1793;
  assign n1795 = G27gat & n1784;
  assign n1796 = ~n1656 & ~n1795;
  assign n1797 = ~G14gat & ~n1796;
  assign n1798 = G14gat & ~n1661;
  assign n1799 = ~n1797 & ~n1798;
  assign n1800 = G21gat & ~n1799;
  assign n1801 = ~n1652 & ~n1800;
  assign n1802 = G8gat & ~n1801;
  assign n1803 = G27gat & n1766;
  assign n1804 = ~G14gat & ~n1803;
  assign n1805 = G14gat & ~n1651;
  assign n1806 = ~n1804 & ~n1805;
  assign n1807 = ~G21gat & ~n1806;
  assign n1808 = G21gat & ~n1774;
  assign n1809 = ~n1807 & ~n1808;
  assign n1810 = ~G8gat & ~n1809;
  assign n1811 = ~n1802 & ~n1810;
  assign n1812 = n171 & ~n1811;
  assign n1813 = ~n1794 & ~n1812;
  assign n1814 = ~G1gat & ~n1813;
  assign n1815 = ~n1764 & ~n1814;
  assign n1816 = G4gat & ~n1815;
  assign n1817 = ~n1696 & ~n1816;
  assign n1818 = keyinput0_G431gat & ~n1817;
  assign n1819 = ~n1348 & ~n1818;
  assign n1820 = keyinput1_G431gat & ~n1819;
  assign n1821 = ~n1347 & ~n1820;
  assign n1822 = keyinput2_G431gat & ~n1821;
  assign n1823 = ~n1344 & ~n1822;
  assign n1824 = keyinput3_G431gat & ~n1823;
  assign G431gat = n1335 | n1824;
  assign n1826 = G11gat & n183;
  assign n1827 = ~keyinput2_G432gat & ~n1826;
  assign n1828 = G37gat & n180;
  assign n1829 = keyinput2_G432gat & ~n1828;
  assign n1830 = ~n1827 & ~n1829;
  assign n1831 = ~keyinput3_G432gat & ~n1830;
  assign n1832 = G63gat & n176;
  assign n1833 = ~keyinput2_G432gat & ~n1832;
  assign n1834 = keyinput2_G432gat & ~n88;
  assign n1835 = ~n1833 & ~n1834;
  assign n1836 = keyinput3_G432gat & ~n1835;
  assign n1837 = ~n1831 & ~n1836;
  assign n1838 = ~keyinput1_G432gat & ~n1837;
  assign n1839 = ~keyinput2_G432gat & ~n137;
  assign n1840 = keyinput2_G432gat & ~n132;
  assign n1841 = ~n1839 & ~n1840;
  assign n1842 = ~keyinput3_G432gat & ~n1841;
  assign n1843 = ~keyinput2_G432gat & n112;
  assign n1844 = G108gat & keyinput2_G432gat;
  assign n1845 = ~n1843 & ~n1844;
  assign n1846 = keyinput3_G432gat & ~n1845;
  assign n1847 = ~n1842 & ~n1846;
  assign n1848 = keyinput1_G432gat & ~n1847;
  assign n1849 = ~n1838 & ~n1848;
  assign n1850 = ~keyinput0_G432gat & ~n1849;
  assign n1851 = keyinput2_G432gat & n865;
  assign n1852 = ~keyinput2_G432gat & ~n867;
  assign n1853 = n868 & n1852;
  assign n1854 = ~n1851 & ~n1853;
  assign n1855 = n160 & ~n1854;
  assign n1856 = ~keyinput3_G432gat & n1855;
  assign n1857 = ~keyinput2_G432gat & ~n133;
  assign n1858 = keyinput2_G432gat & n72;
  assign n1859 = ~n1857 & ~n1858;
  assign n1860 = keyinput3_G432gat & ~n1859;
  assign n1861 = ~n1856 & ~n1860;
  assign n1862 = ~keyinput1_G432gat & ~n1861;
  assign n1863 = ~keyinput2_G432gat & ~n181;
  assign n1864 = keyinput2_G432gat & n160;
  assign n1865 = ~n1863 & ~n1864;
  assign n1866 = ~keyinput3_G432gat & ~n1865;
  assign n1867 = ~keyinput2_G432gat & ~n111;
  assign n1868 = n430 & ~n477;
  assign n1869 = n524 & ~n571;
  assign n1870 = ~n1868 & ~n1869;
  assign n1871 = ~n618 & n1870;
  assign n1872 = G40gat & ~n1871;
  assign n1873 = ~G34gat & n1872;
  assign n1874 = ~G66gat & n1868;
  assign n1875 = n92 & n173;
  assign n1876 = ~n281 & n1875;
  assign n1877 = G92gat & n430;
  assign n1878 = n281 & n1877;
  assign n1879 = ~n1876 & ~n1878;
  assign n1880 = ~n524 & n1879;
  assign n1881 = G66gat & ~n1880;
  assign n1882 = ~n1874 & ~n1881;
  assign n1883 = n311 & n1882;
  assign n1884 = ~n1355 & n1879;
  assign n1885 = n74 & ~n430;
  assign n1886 = ~n477 & ~n1885;
  assign n1887 = G79gat & ~n1886;
  assign n1888 = n295 & n1887;
  assign n1889 = ~n1884 & ~n1888;
  assign n1890 = ~n311 & ~n1889;
  assign n1891 = ~n1883 & ~n1890;
  assign n1892 = ~n327 & ~n1891;
  assign n1893 = ~n524 & ~n1886;
  assign n1894 = n571 & ~n1868;
  assign n1895 = ~n1893 & ~n1894;
  assign n1896 = G53gat & ~n1895;
  assign n1897 = n327 & n1896;
  assign n1898 = ~n1892 & ~n1897;
  assign n1899 = ~G40gat & n1898;
  assign n1900 = n173 & n216;
  assign n1901 = n73 & ~n1900;
  assign n1902 = ~n281 & ~n1901;
  assign n1903 = ~n1877 & ~n1902;
  assign n1904 = ~G79gat & ~n1903;
  assign n1905 = ~G73gat & ~n1887;
  assign n1906 = ~G86gat & n1877;
  assign n1907 = ~G92gat & n1875;
  assign n1908 = G86gat & n1907;
  assign n1909 = ~n1906 & ~n1908;
  assign n1910 = ~G76gat & ~n1909;
  assign n1911 = G82gat & n1910;
  assign n1912 = ~n78 & ~n92;
  assign n1913 = n173 & ~n1912;
  assign n1914 = ~n895 & n1913;
  assign n1915 = ~n1911 & ~n1914;
  assign n1916 = ~n908 & ~n1915;
  assign n1917 = ~n1905 & ~n1916;
  assign n1918 = ~n1904 & n1917;
  assign n1919 = ~n177 & n1915;
  assign n1920 = ~n1918 & ~n1919;
  assign n1921 = ~n178 & n1920;
  assign n1922 = ~G60gat & ~n1882;
  assign n1923 = ~n295 & n1915;
  assign n1924 = ~n1888 & ~n1923;
  assign n1925 = ~G66gat & n1924;
  assign n1926 = G66gat & n1920;
  assign n1927 = ~n1925 & ~n1926;
  assign n1928 = G60gat & ~n1927;
  assign n1929 = ~n1922 & ~n1928;
  assign n1930 = n178 & ~n1929;
  assign n1931 = ~n1921 & ~n1930;
  assign n1932 = ~n903 & n1931;
  assign n1933 = ~G47gat & n1896;
  assign n1934 = ~n295 & n1903;
  assign n1935 = ~n1888 & ~n1934;
  assign n1936 = ~n311 & n1935;
  assign n1937 = ~G50gat & n1922;
  assign n1938 = G56gat & n1937;
  assign n1939 = ~n1936 & ~n1938;
  assign n1940 = ~G53gat & n1939;
  assign n1941 = G47gat & n1940;
  assign n1942 = ~n1933 & ~n1941;
  assign n1943 = n172 & ~n1942;
  assign n1944 = ~n1932 & ~n1943;
  assign n1945 = G40gat & n1944;
  assign n1946 = ~n1899 & ~n1945;
  assign n1947 = G34gat & ~n1946;
  assign n1948 = ~n1873 & ~n1947;
  assign n1949 = ~G24gat & ~n1948;
  assign n1950 = G95gat & n99;
  assign n1951 = ~n174 & n1950;
  assign n1952 = G92gat & n1913;
  assign n1953 = ~n1907 & ~n1952;
  assign n1954 = G86gat & ~n1953;
  assign n1955 = ~n1906 & ~n1954;
  assign n1956 = ~G76gat & ~n1955;
  assign n1957 = G82gat & n1956;
  assign n1958 = ~n1951 & ~n1957;
  assign n1959 = ~G69gat & ~n1958;
  assign n1960 = ~n94 & ~n173;
  assign n1961 = ~n1950 & ~n1960;
  assign n1962 = ~G76gat & ~n865;
  assign n1963 = G82gat & n1962;
  assign n1964 = ~n1961 & ~n1963;
  assign n1965 = ~n1911 & ~n1964;
  assign n1966 = G79gat & ~n1965;
  assign n1967 = ~n1904 & ~n1966;
  assign n1968 = G73gat & ~n1967;
  assign n1969 = ~n1905 & ~n1968;
  assign n1970 = ~G63gat & ~n1969;
  assign n1971 = G63gat & ~n1958;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = G69gat & ~n1972;
  assign n1974 = ~n1959 & ~n1973;
  assign n1975 = ~n178 & ~n1974;
  assign n1976 = ~n177 & n1958;
  assign n1977 = G79gat & ~n1958;
  assign n1978 = ~n1904 & ~n1977;
  assign n1979 = G73gat & ~n1978;
  assign n1980 = ~n1905 & ~n1979;
  assign n1981 = n177 & n1980;
  assign n1982 = ~n1976 & ~n1981;
  assign n1983 = G66gat & n1982;
  assign n1984 = ~n1925 & ~n1983;
  assign n1985 = G60gat & ~n1984;
  assign n1986 = ~n1922 & ~n1985;
  assign n1987 = ~G50gat & ~n1986;
  assign n1988 = G56gat & n1987;
  assign n1989 = ~n1975 & ~n1988;
  assign n1990 = ~n172 & ~n1989;
  assign n1991 = ~n177 & ~n1965;
  assign n1992 = G69gat & n1970;
  assign n1993 = ~n1991 & ~n1992;
  assign n1994 = ~n178 & n1993;
  assign n1995 = G66gat & ~n1993;
  assign n1996 = ~n1925 & ~n1995;
  assign n1997 = G60gat & ~n1996;
  assign n1998 = ~n1922 & ~n1997;
  assign n1999 = n178 & n1998;
  assign n2000 = ~n1994 & ~n1999;
  assign n2001 = G53gat & ~n2000;
  assign n2002 = ~n1940 & ~n2001;
  assign n2003 = G47gat & ~n2002;
  assign n2004 = ~n1933 & ~n2003;
  assign n2005 = ~G37gat & n2004;
  assign n2006 = G43gat & n2005;
  assign n2007 = ~n1990 & ~n2006;
  assign n2008 = ~G40gat & ~n2007;
  assign n2009 = ~G92gat & n1950;
  assign n2010 = n1509 & n2009;
  assign n2011 = ~n1956 & ~n2010;
  assign n2012 = G82gat & ~n2011;
  assign n2013 = n202 & n243;
  assign n2014 = ~n99 & ~n2013;
  assign n2015 = G95gat & ~n2014;
  assign n2016 = ~n815 & n2015;
  assign n2017 = ~n2012 & ~n2016;
  assign n2018 = ~G69gat & ~n2017;
  assign n2019 = ~n270 & ~n1950;
  assign n2020 = ~n174 & ~n2019;
  assign n2021 = ~n1957 & ~n2020;
  assign n2022 = ~G79gat & ~n2021;
  assign n2023 = ~G73gat & n2022;
  assign n2024 = ~n523 & ~n2017;
  assign n2025 = ~n2023 & ~n2024;
  assign n2026 = G63gat & ~n2025;
  assign n2027 = ~n1970 & ~n2026;
  assign n2028 = G69gat & ~n2027;
  assign n2029 = ~n2018 & ~n2028;
  assign n2030 = ~G56gat & ~n2029;
  assign n2031 = ~n820 & ~n2029;
  assign n2032 = ~n177 & ~n2017;
  assign n2033 = ~n1992 & ~n2032;
  assign n2034 = ~G66gat & ~n2033;
  assign n2035 = ~G60gat & n2034;
  assign n2036 = ~n2031 & ~n2035;
  assign n2037 = G50gat & ~n2036;
  assign n2038 = ~n1987 & ~n2037;
  assign n2039 = G56gat & ~n2038;
  assign n2040 = ~n2030 & ~n2039;
  assign n2041 = ~G43gat & ~n2040;
  assign n2042 = ~n617 & n2040;
  assign n2043 = ~n177 & ~n2021;
  assign n2044 = ~n1992 & ~n2043;
  assign n2045 = ~n178 & ~n2044;
  assign n2046 = ~n1988 & ~n2045;
  assign n2047 = n617 & n2046;
  assign n2048 = ~n2042 & ~n2047;
  assign n2049 = G37gat & n2048;
  assign n2050 = ~n2005 & ~n2049;
  assign n2051 = G43gat & ~n2050;
  assign n2052 = ~n2041 & ~n2051;
  assign n2053 = G40gat & ~n2052;
  assign n2054 = ~n2008 & ~n2053;
  assign n2055 = ~G34gat & ~n2054;
  assign n2056 = G89gat & n106;
  assign n2057 = ~n99 & ~n2056;
  assign n2058 = G95gat & ~n2057;
  assign n2059 = ~G82gat & n2058;
  assign n2060 = G92gat & n2015;
  assign n2061 = ~n2009 & ~n2060;
  assign n2062 = ~G86gat & ~n2061;
  assign n2063 = G86gat & n2058;
  assign n2064 = ~n2062 & ~n2063;
  assign n2065 = G76gat & ~n2064;
  assign n2066 = ~n1956 & ~n2065;
  assign n2067 = G82gat & ~n2066;
  assign n2068 = ~n2059 & ~n2067;
  assign n2069 = ~G69gat & ~n2068;
  assign n2070 = ~G95gat & ~n103;
  assign n2071 = G99gat & ~n103;
  assign n2072 = ~n106 & ~n2071;
  assign n2073 = G89gat & ~n2072;
  assign n2074 = ~n99 & ~n2073;
  assign n2075 = G95gat & ~n2074;
  assign n2076 = ~n2070 & ~n2075;
  assign n2077 = ~G82gat & ~n2076;
  assign n2078 = ~n476 & n2076;
  assign n2079 = n476 & ~n1950;
  assign n2080 = ~n2078 & ~n2079;
  assign n2081 = G76gat & n2080;
  assign n2082 = ~n1956 & ~n2081;
  assign n2083 = G82gat & ~n2082;
  assign n2084 = ~n2077 & ~n2083;
  assign n2085 = G79gat & ~n2084;
  assign n2086 = ~n2022 & ~n2085;
  assign n2087 = ~G73gat & ~n2086;
  assign n2088 = G73gat & ~n2068;
  assign n2089 = ~n2087 & ~n2088;
  assign n2090 = G63gat & ~n2089;
  assign n2091 = ~n1970 & ~n2090;
  assign n2092 = G69gat & ~n2091;
  assign n2093 = ~n2069 & ~n2092;
  assign n2094 = ~G56gat & ~n2093;
  assign n2095 = ~n523 & ~n2068;
  assign n2096 = ~n2023 & ~n2095;
  assign n2097 = G63gat & ~n2096;
  assign n2098 = ~n1970 & ~n2097;
  assign n2099 = G69gat & ~n2098;
  assign n2100 = ~n2069 & ~n2099;
  assign n2101 = G66gat & ~n2100;
  assign n2102 = ~n2034 & ~n2101;
  assign n2103 = ~G60gat & ~n2102;
  assign n2104 = G60gat & ~n2093;
  assign n2105 = ~n2103 & ~n2104;
  assign n2106 = G50gat & ~n2105;
  assign n2107 = ~n1987 & ~n2106;
  assign n2108 = G56gat & ~n2107;
  assign n2109 = ~n2094 & ~n2108;
  assign n2110 = ~G43gat & ~n2109;
  assign n2111 = ~G53gat & ~n2046;
  assign n2112 = ~G69gat & ~n2084;
  assign n2113 = G73gat & ~n2084;
  assign n2114 = ~n2087 & ~n2113;
  assign n2115 = G63gat & ~n2114;
  assign n2116 = ~n1970 & ~n2115;
  assign n2117 = G69gat & ~n2116;
  assign n2118 = ~n2112 & ~n2117;
  assign n2119 = ~G56gat & ~n2118;
  assign n2120 = ~n820 & ~n2118;
  assign n2121 = ~n2035 & ~n2120;
  assign n2122 = G50gat & ~n2121;
  assign n2123 = ~n1987 & ~n2122;
  assign n2124 = G56gat & ~n2123;
  assign n2125 = ~n2119 & ~n2124;
  assign n2126 = G53gat & ~n2125;
  assign n2127 = ~n2111 & ~n2126;
  assign n2128 = ~G47gat & ~n2127;
  assign n2129 = G47gat & ~n2109;
  assign n2130 = ~n2128 & ~n2129;
  assign n2131 = G37gat & ~n2130;
  assign n2132 = ~n2005 & ~n2131;
  assign n2133 = G43gat & ~n2132;
  assign n2134 = ~n2110 & ~n2133;
  assign n2135 = ~G40gat & ~n2134;
  assign n2136 = ~n99 & ~n109;
  assign n2137 = G95gat & ~n2136;
  assign n2138 = ~G82gat & n2137;
  assign n2139 = ~G92gat & n2058;
  assign n2140 = G92gat & n2137;
  assign n2141 = ~n2139 & ~n2140;
  assign n2142 = G86gat & ~n2141;
  assign n2143 = ~n2062 & ~n2142;
  assign n2144 = G76gat & ~n2143;
  assign n2145 = ~n1956 & ~n2144;
  assign n2146 = G82gat & ~n2145;
  assign n2147 = ~n2138 & ~n2146;
  assign n2148 = ~G69gat & ~n2147;
  assign n2149 = ~G95gat & ~n88;
  assign n2150 = ~n89 & ~n106;
  assign n2151 = G89gat & ~n2150;
  assign n2152 = ~n99 & ~n2151;
  assign n2153 = G95gat & ~n2152;
  assign n2154 = ~n2149 & ~n2153;
  assign n2155 = ~G82gat & ~n2154;
  assign n2156 = G86gat & ~n2154;
  assign n2157 = ~n2062 & ~n2156;
  assign n2158 = G76gat & ~n2157;
  assign n2159 = ~n1956 & ~n2158;
  assign n2160 = G82gat & ~n2159;
  assign n2161 = ~n2155 & ~n2160;
  assign n2162 = ~G79gat & ~n2161;
  assign n2163 = G79gat & ~n2147;
  assign n2164 = ~n2162 & ~n2163;
  assign n2165 = G73gat & ~n2164;
  assign n2166 = ~n2087 & ~n2165;
  assign n2167 = G63gat & ~n2166;
  assign n2168 = ~n1970 & ~n2167;
  assign n2169 = G69gat & ~n2168;
  assign n2170 = ~n2148 & ~n2169;
  assign n2171 = ~G56gat & ~n2170;
  assign n2172 = G73gat & ~n2147;
  assign n2173 = ~n2087 & ~n2172;
  assign n2174 = G63gat & ~n2173;
  assign n2175 = ~n1970 & ~n2174;
  assign n2176 = G69gat & ~n2175;
  assign n2177 = ~n2148 & ~n2176;
  assign n2178 = ~G66gat & ~n2177;
  assign n2179 = G66gat & ~n2170;
  assign n2180 = ~n2178 & ~n2179;
  assign n2181 = G60gat & ~n2180;
  assign n2182 = ~n2103 & ~n2181;
  assign n2183 = G50gat & ~n2182;
  assign n2184 = ~n1987 & ~n2183;
  assign n2185 = G56gat & ~n2184;
  assign n2186 = ~n2171 & ~n2185;
  assign n2187 = ~G43gat & ~n2186;
  assign n2188 = ~G69gat & ~n2161;
  assign n2189 = G73gat & ~n2161;
  assign n2190 = ~n2087 & ~n2189;
  assign n2191 = G63gat & ~n2190;
  assign n2192 = ~n1970 & ~n2191;
  assign n2193 = G69gat & ~n2192;
  assign n2194 = ~n2188 & ~n2193;
  assign n2195 = ~G56gat & ~n2194;
  assign n2196 = G60gat & ~n2194;
  assign n2197 = ~n2103 & ~n2196;
  assign n2198 = G50gat & ~n2197;
  assign n2199 = ~n1987 & ~n2198;
  assign n2200 = G56gat & ~n2199;
  assign n2201 = ~n2195 & ~n2200;
  assign n2202 = ~G53gat & ~n2201;
  assign n2203 = G53gat & ~n2186;
  assign n2204 = ~n2202 & ~n2203;
  assign n2205 = G47gat & ~n2204;
  assign n2206 = ~n2128 & ~n2205;
  assign n2207 = G37gat & ~n2206;
  assign n2208 = ~n2005 & ~n2207;
  assign n2209 = G43gat & ~n2208;
  assign n2210 = ~n2187 & ~n2209;
  assign n2211 = G40gat & ~n2210;
  assign n2212 = ~n2135 & ~n2211;
  assign n2213 = G34gat & ~n2212;
  assign n2214 = ~n2055 & ~n2213;
  assign n2215 = G24gat & ~n2214;
  assign n2216 = ~n1949 & ~n2215;
  assign n2217 = G30gat & ~n2216;
  assign n2218 = ~G95gat & ~n111;
  assign n2219 = G95gat & ~n116;
  assign n2220 = ~n2218 & ~n2219;
  assign n2221 = ~G82gat & ~n2220;
  assign n2222 = G92gat & ~n2220;
  assign n2223 = ~n2139 & ~n2222;
  assign n2224 = G86gat & ~n2223;
  assign n2225 = ~n2062 & ~n2224;
  assign n2226 = G76gat & ~n2225;
  assign n2227 = ~n1956 & ~n2226;
  assign n2228 = G82gat & ~n2227;
  assign n2229 = ~n2221 & ~n2228;
  assign n2230 = ~G69gat & ~n2229;
  assign n2231 = G79gat & ~n2229;
  assign n2232 = ~n2162 & ~n2231;
  assign n2233 = G73gat & ~n2232;
  assign n2234 = ~n2087 & ~n2233;
  assign n2235 = G63gat & ~n2234;
  assign n2236 = ~n1970 & ~n2235;
  assign n2237 = G69gat & ~n2236;
  assign n2238 = ~n2230 & ~n2237;
  assign n2239 = ~G56gat & ~n2238;
  assign n2240 = G66gat & ~n2238;
  assign n2241 = ~n2178 & ~n2240;
  assign n2242 = G60gat & ~n2241;
  assign n2243 = ~n2103 & ~n2242;
  assign n2244 = G50gat & ~n2243;
  assign n2245 = ~n1987 & ~n2244;
  assign n2246 = G56gat & ~n2245;
  assign n2247 = ~n2239 & ~n2246;
  assign n2248 = G53gat & ~n2247;
  assign n2249 = ~n2202 & ~n2248;
  assign n2250 = G47gat & ~n2249;
  assign n2251 = ~n2128 & ~n2250;
  assign n2252 = G37gat & ~n2251;
  assign n2253 = ~n2005 & ~n2252;
  assign n2254 = G43gat & ~n2253;
  assign n2255 = ~G82gat & n2219;
  assign n2256 = ~n2146 & ~n2255;
  assign n2257 = ~G69gat & ~n2256;
  assign n2258 = ~n2237 & ~n2257;
  assign n2259 = ~G56gat & ~n2258;
  assign n2260 = ~n870 & ~n2256;
  assign n2261 = G73gat & n2162;
  assign n2262 = ~n2087 & ~n2261;
  assign n2263 = G63gat & ~n2262;
  assign n2264 = ~n1970 & ~n2263;
  assign n2265 = G69gat & ~n2264;
  assign n2266 = ~n2260 & ~n2265;
  assign n2267 = G66gat & ~n2266;
  assign n2268 = ~n2178 & ~n2267;
  assign n2269 = G60gat & ~n2268;
  assign n2270 = ~n2103 & ~n2269;
  assign n2271 = G50gat & ~n2270;
  assign n2272 = ~n1987 & ~n2271;
  assign n2273 = G56gat & ~n2272;
  assign n2274 = ~n2259 & ~n2273;
  assign n2275 = ~G43gat & ~n2274;
  assign n2276 = ~n2254 & ~n2275;
  assign n2277 = ~G30gat & ~n2276;
  assign n2278 = ~n2217 & ~n2277;
  assign n2279 = ~G17gat & ~n2278;
  assign n2280 = ~n618 & ~n1895;
  assign n2281 = ~n665 & ~n2280;
  assign n2282 = G27gat & ~n2281;
  assign n2283 = ~G21gat & ~n2282;
  assign n2284 = ~n1157 & ~n1939;
  assign n2285 = n1157 & ~n1896;
  assign n2286 = ~n2284 & ~n2285;
  assign n2287 = ~n343 & ~n2286;
  assign n2288 = n343 & n1872;
  assign n2289 = ~n2287 & ~n2288;
  assign n2290 = ~G27gat & ~n2289;
  assign n2291 = ~n903 & ~n2000;
  assign n2292 = ~n1943 & ~n2291;
  assign n2293 = ~n897 & n2292;
  assign n2294 = G34gat & n1899;
  assign n2295 = ~n1873 & ~n2294;
  assign n2296 = n182 & ~n2295;
  assign n2297 = ~n2293 & ~n2296;
  assign n2298 = G27gat & ~n2297;
  assign n2299 = ~n2290 & ~n2298;
  assign n2300 = G21gat & ~n2299;
  assign n2301 = ~n2283 & ~n2300;
  assign n2302 = ~G11gat & ~n2301;
  assign n2303 = ~n172 & n2046;
  assign n2304 = n172 & ~n2004;
  assign n2305 = ~n2303 & ~n2304;
  assign n2306 = ~n182 & ~n2305;
  assign n2307 = ~G24gat & n1948;
  assign n2308 = G30gat & n2307;
  assign n2309 = ~n2306 & ~n2308;
  assign n2310 = ~G27gat & n2309;
  assign n2311 = ~G40gat & n2007;
  assign n2312 = n1697 & n2311;
  assign n2313 = ~n2307 & ~n2312;
  assign n2314 = G30gat & ~n2313;
  assign n2315 = G47gat & ~n2125;
  assign n2316 = ~n2128 & ~n2315;
  assign n2317 = G37gat & ~n2316;
  assign n2318 = ~n2005 & ~n2317;
  assign n2319 = G43gat & n2318;
  assign n2320 = ~G43gat & n2125;
  assign n2321 = ~n2319 & ~n2320;
  assign n2322 = ~n826 & ~n2321;
  assign n2323 = ~n2314 & ~n2322;
  assign n2324 = G27gat & n2323;
  assign n2325 = ~n2310 & ~n2324;
  assign n2326 = ~G21gat & ~n2325;
  assign n2327 = n1697 & n2054;
  assign n2328 = ~n2307 & ~n2327;
  assign n2329 = G30gat & ~n2328;
  assign n2330 = ~G43gat & n2201;
  assign n2331 = G47gat & ~n2201;
  assign n2332 = ~n2128 & ~n2331;
  assign n2333 = G37gat & ~n2332;
  assign n2334 = ~n2005 & ~n2333;
  assign n2335 = G43gat & n2334;
  assign n2336 = ~n2330 & ~n2335;
  assign n2337 = ~n845 & ~n2336;
  assign n2338 = ~G27gat & ~n2337;
  assign n2339 = ~n2329 & n2338;
  assign n2340 = ~G43gat & ~n2247;
  assign n2341 = ~n2254 & ~n2340;
  assign n2342 = ~n861 & ~n2341;
  assign n2343 = G34gat & n2135;
  assign n2344 = ~n2055 & ~n2343;
  assign n2345 = G24gat & ~n2344;
  assign n2346 = ~n1949 & ~n2345;
  assign n2347 = G30gat & ~n2346;
  assign n2348 = ~n2342 & ~n2347;
  assign n2349 = G27gat & ~n2348;
  assign n2350 = ~n2339 & ~n2349;
  assign n2351 = G21gat & ~n2350;
  assign n2352 = ~n2326 & ~n2351;
  assign n2353 = G11gat & ~n2352;
  assign n2354 = ~n2302 & ~n2353;
  assign n2355 = G17gat & ~n2354;
  assign n2356 = ~n2279 & ~n2355;
  assign n2357 = ~G4gat & ~n2356;
  assign n2358 = ~n897 & n1944;
  assign n2359 = ~n2296 & ~n2358;
  assign n2360 = ~G14gat & n2359;
  assign n2361 = ~n182 & ~n2007;
  assign n2362 = G30gat & n1949;
  assign n2363 = ~n2361 & ~n2362;
  assign n2364 = G14gat & n2363;
  assign n2365 = ~n2360 & ~n2364;
  assign n2366 = G8gat & ~n2365;
  assign n2367 = ~n665 & ~n1871;
  assign n2368 = ~G14gat & n2367;
  assign n2369 = ~n343 & n1898;
  assign n2370 = ~n2288 & ~n2369;
  assign n2371 = G14gat & ~n2370;
  assign n2372 = ~n2368 & ~n2371;
  assign n2373 = ~G8gat & n2372;
  assign n2374 = ~n2366 & ~n2373;
  assign n2375 = ~n171 & ~n2374;
  assign n2376 = G27gat & ~n2359;
  assign n2377 = ~n2290 & ~n2376;
  assign n2378 = ~G14gat & ~n2377;
  assign n2379 = G14gat & ~n2299;
  assign n2380 = ~n2378 & ~n2379;
  assign n2381 = G21gat & ~n2380;
  assign n2382 = ~n2283 & ~n2381;
  assign n2383 = G8gat & n2382;
  assign n2384 = G27gat & ~n2368;
  assign n2385 = G14gat & n2281;
  assign n2386 = n2384 & ~n2385;
  assign n2387 = ~G21gat & ~n2386;
  assign n2388 = G21gat & ~n2372;
  assign n2389 = ~n2387 & ~n2388;
  assign n2390 = ~G8gat & n2389;
  assign n2391 = ~n2383 & ~n2390;
  assign n2392 = n171 & ~n2391;
  assign n2393 = ~n2375 & ~n2392;
  assign n2394 = ~G1gat & n2393;
  assign n2395 = n1697 & n2008;
  assign n2396 = ~n1949 & ~n2395;
  assign n2397 = G30gat & ~n2396;
  assign n2398 = ~n826 & ~n2052;
  assign n2399 = ~n2397 & ~n2398;
  assign n2400 = ~G14gat & ~n2399;
  assign n2401 = ~G30gat & ~n2134;
  assign n2402 = G34gat & ~n2134;
  assign n2403 = ~n2055 & ~n2402;
  assign n2404 = G24gat & ~n2403;
  assign n2405 = ~n1949 & ~n2404;
  assign n2406 = G30gat & ~n2405;
  assign n2407 = ~n2401 & ~n2406;
  assign n2408 = G14gat & ~n2407;
  assign n2409 = ~n2400 & ~n2408;
  assign n2410 = ~G8gat & ~n2409;
  assign n2411 = ~G30gat & ~n2210;
  assign n2412 = ~n2217 & ~n2411;
  assign n2413 = ~G14gat & ~n2412;
  assign n2414 = G14gat & ~n2278;
  assign n2415 = ~n2413 & ~n2414;
  assign n2416 = G8gat & ~n2415;
  assign n2417 = ~n2410 & ~n2416;
  assign n2418 = ~G17gat & ~n2417;
  assign n2419 = G27gat & ~n2399;
  assign n2420 = ~n2310 & ~n2419;
  assign n2421 = ~G14gat & ~n2420;
  assign n2422 = G14gat & ~n2325;
  assign n2423 = ~n2421 & ~n2422;
  assign n2424 = ~G21gat & ~n2423;
  assign n2425 = G21gat & ~n2409;
  assign n2426 = ~n2424 & ~n2425;
  assign n2427 = ~G8gat & ~n2426;
  assign n2428 = G14gat & ~n2348;
  assign n2429 = ~n2413 & ~n2428;
  assign n2430 = G27gat & ~n2429;
  assign n2431 = ~n2339 & ~n2430;
  assign n2432 = G21gat & ~n2431;
  assign n2433 = ~n2326 & ~n2432;
  assign n2434 = G8gat & ~n2433;
  assign n2435 = ~n2427 & ~n2434;
  assign n2436 = G11gat & ~n2435;
  assign n2437 = ~n2302 & ~n2436;
  assign n2438 = G17gat & ~n2437;
  assign n2439 = ~n2418 & ~n2438;
  assign n2440 = G1gat & ~n2439;
  assign n2441 = ~n2394 & ~n2440;
  assign n2442 = G4gat & ~n2441;
  assign n2443 = ~n2357 & ~n2442;
  assign n2444 = keyinput2_G432gat & ~n2443;
  assign n2445 = ~n1867 & ~n2444;
  assign n2446 = keyinput3_G432gat & ~n2445;
  assign n2447 = ~n1866 & ~n2446;
  assign n2448 = keyinput1_G432gat & ~n2447;
  assign n2449 = ~n1862 & ~n2448;
  assign n2450 = keyinput0_G432gat & ~n2449;
  assign G432gat = n1850 | n2450;
endmodule


