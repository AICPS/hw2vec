// Verilog File 
module top (G1gat,G8gat,G13gat,G17gat,G26gat,G29gat,G36gat,G42gat,G51gat,
G55gat,G59gat,G68gat,G72gat,G73gat,G74gat,G75gat,G80gat,G85gat,G86gat,
G87gat,G88gat,G89gat,G90gat,G91gat,G96gat,G101gat,G106gat,G111gat,G116gat,
G121gat,G126gat,G130gat,G135gat,G138gat,G143gat,G146gat,G149gat,G152gat,G153gat,
G156gat,G159gat,G165gat,G171gat,G177gat,G183gat,G189gat,G195gat,G201gat,G207gat,
G210gat,G219gat,G228gat,G237gat,G246gat,G255gat,G259gat,G260gat,G261gat,G267gat,
G268gat,G388gat,G389gat,G390gat,G391gat,G418gat,G419gat,G420gat,G421gat,G422gat,
G423gat,G446gat,G447gat,G448gat,G449gat,G450gat,G767gat,G768gat,G850gat,G863gat,
G864gat,G865gat,G866gat,G874gat,G878gat,G879gat,G880gat,keyinput0,keyinput1,keyinput2,
keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,
keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,
keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,
keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,
keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,
keyinput53,keyinput54,keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,
keyinput63,keyinput64,keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,
keyinput73,keyinput74,keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,
keyinput83,keyinput84,keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,
keyinput93,keyinput94,keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,
keyinput103,keyinput104,keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,
keyinput113,keyinput114,keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,
keyinput123,keyinput124,keyinput125,keyinput126,keyinput127,keyinput128,keyinput129,keyinput130,keyinput131,keyinput132,
keyinput133,keyinput134,keyinput135,keyinput136,keyinput137,keyinput138,keyinput139,keyinput140,keyinput141,keyinput142,
keyinput143,keyinput144,keyinput145,keyinput146,keyinput147,keyinput148,keyinput149,keyinput150,keyinput151,keyinput152,
keyinput153,keyinput154,keyinput155,keyinput156,keyinput157,keyinput158,keyinput159,keyinput160,keyinput161,keyinput162,
keyinput163,keyinput164,keyinput165,keyinput166,keyinput167,keyinput168,keyinput169,keyinput170,keyinput171,keyinput172,
keyinput173,keyinput174,keyinput175,keyinput176,keyinput177,keyinput178,keyinput179,keyinput180,keyinput181,keyinput182,
keyinput183,keyinput184,keyinput185,keyinput186,keyinput187,keyinput188,keyinput189,keyinput190,keyinput191,keyinput192,
keyinput193,keyinput194,keyinput195,keyinput196,keyinput197,keyinput198,keyinput199,keyinput200,keyinput201,keyinput202);

input G1gat,G8gat,G13gat,G17gat,G26gat,G29gat,G36gat,G42gat,G51gat,
G55gat,G59gat,G68gat,G72gat,G73gat,G74gat,G75gat,G80gat,G85gat,G86gat,
G87gat,G88gat,G89gat,G90gat,G91gat,G96gat,G101gat,G106gat,G111gat,G116gat,
G121gat,G126gat,G130gat,G135gat,G138gat,G143gat,G146gat,G149gat,G152gat,G153gat,
G156gat,G159gat,G165gat,G171gat,G177gat,G183gat,G189gat,G195gat,G201gat,G207gat,
G210gat,G219gat,G228gat,G237gat,G246gat,G255gat,G259gat,G260gat,G261gat,G267gat,
G268gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,
keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,
keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,
keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,keyinput38,
keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,keyinput48,
keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,keyinput55,keyinput56,keyinput57,keyinput58,
keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,keyinput65,keyinput66,keyinput67,keyinput68,
keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,keyinput75,keyinput76,keyinput77,keyinput78,
keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,keyinput85,keyinput86,keyinput87,keyinput88,
keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,keyinput95,keyinput96,keyinput97,keyinput98,
keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,keyinput105,keyinput106,keyinput107,keyinput108,
keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,keyinput115,keyinput116,keyinput117,keyinput118,
keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,keyinput125,keyinput126,keyinput127,keyinput128,
keyinput129,keyinput130,keyinput131,keyinput132,keyinput133,keyinput134,keyinput135,keyinput136,keyinput137,keyinput138,
keyinput139,keyinput140,keyinput141,keyinput142,keyinput143,keyinput144,keyinput145,keyinput146,keyinput147,keyinput148,
keyinput149,keyinput150,keyinput151,keyinput152,keyinput153,keyinput154,keyinput155,keyinput156,keyinput157,keyinput158,
keyinput159,keyinput160,keyinput161,keyinput162,keyinput163,keyinput164,keyinput165,keyinput166,keyinput167,keyinput168,
keyinput169,keyinput170,keyinput171,keyinput172,keyinput173,keyinput174,keyinput175,keyinput176,keyinput177,keyinput178,
keyinput179,keyinput180,keyinput181,keyinput182,keyinput183,keyinput184,keyinput185,keyinput186,keyinput187,keyinput188,
keyinput189,keyinput190,keyinput191,keyinput192,keyinput193,keyinput194,keyinput195,keyinput196,keyinput197,keyinput198,
keyinput199,keyinput200,keyinput201,keyinput202;

output G388gat,G389gat,G390gat,G391gat,G418gat,G419gat,G420gat,G421gat,G422gat,
G423gat,G446gat,G447gat,G448gat,G449gat,G450gat,G767gat,G768gat,G850gat,G863gat,
G864gat,G865gat,G866gat,G874gat,G878gat,G879gat,G880gat;

wire G269gat,G270gat,G273gat,G276gat,G279gat,G280gat,G284gat,G285gat,G286gat,
G287gat,G290gat,G291gat,G292gat,G293gat,G294gat,G295gat,G296gat,G297gat,G298gat,
G301gat,G302gat,G303gat,G304gat,G305gat,G306gat,G307gat,G308gat,G309gat,G310gat,
G316gat,G317gat,G318gat,G319gat,G322gat,G323gat,G324gat,G325gat,G326gat,G327gat,
G328gat,G329gat,G330gat,G331gat,G332gat,G333gat,G334gat,G335gat,G336gat,G337gat,
G338gat,G339gat,G340gat,G341gat,G342gat,G343gat,G344gat,G345gat,G346gat,G347gat,
G348gat,G349gat,G350gat,G351gat,G352gat,G353gat,G354gat,G355gat,G356gat,G357gat,
G360gat,G363gat,G366gat,G369gat,G375gat,G376gat,G379gat,G382gat,G385gat,G392gat,
G393gat,G399gat,G400gat,G401gat,G402gat,G403gat,G404gat,G405gat,G406gat,G407gat,
G408gat,G409gat,G410gat,G411gat,G412gat,G413gat,G414gat,G415gat,G416gat,G417gat,
G424gat,G425gat,G426gat,G427gat,G432gat,G437gat,G442gat,G443gat,G444gat,G445gat,
G451gat,G460gat,G463gat,G466gat,G475gat,G476gat,G477gat,G478gat,G479gat,G480gat,
G481gat,G482gat,G483gat,G488gat,G489gat,G490gat,G491gat,G492gat,G495gat,G498gat,
G499gat,G500gat,G501gat,G502gat,G503gat,G504gat,G505gat,G506gat,G507gat,G508gat,
G509gat,G510gat,G511gat,G512gat,G513gat,G514gat,G515gat,G516gat,G517gat,G518gat,
G519gat,G520gat,G521gat,G522gat,G523gat,G524gat,G525gat,G526gat,G527gat,G528gat,
G529gat,G530gat,G533gat,G536gat,G537gat,G538gat,G539gat,G540gat,G541gat,G542gat,
G543gat,G544gat,G547gat,G550gat,G551gat,G552gat,G553gat,G557gat,G561gat,G565gat,
G569gat,G573gat,G577gat,G581gat,G585gat,G586gat,G587gat,G588gat,G589gat,G590gat,
G593gat,G596gat,G597gat,G600gat,G605gat,G606gat,G609gat,G615gat,G616gat,G619gat,
G624gat,G625gat,G628gat,G631gat,G632gat,G635gat,G640gat,G641gat,G644gat,G650gat,
G651gat,G654gat,G659gat,G660gat,G661gat,G662gat,G665gat,G669gat,G670gat,G673gat,
G677gat,G678gat,G682gat,G686gat,G687gat,G692gat,G696gat,G697gat,G700gat,G704gat,
G705gat,G708gat,G712gat,G713gat,G717gat,G721gat,G722gat,G727gat,G731gat,G732gat,
G733gat,G734gat,G735gat,G736gat,G737gat,G738gat,G739gat,G740gat,G741gat,G742gat,
G743gat,G744gat,G745gat,G746gat,G747gat,G748gat,G749gat,G750gat,G751gat,G752gat,
G753gat,G754gat,G755gat,G756gat,G757gat,G758gat,G759gat,G760gat,G761gat,G762gat,
G763gat,G764gat,G765gat,G766gat,G769gat,G770gat,G771gat,G772gat,G773gat,G777gat,
G778gat,G781gat,G782gat,G785gat,G786gat,G787gat,G788gat,G789gat,G790gat,G791gat,
G792gat,G793gat,G794gat,G795gat,G796gat,G802gat,G803gat,G804gat,G805gat,G806gat,
G807gat,G808gat,G809gat,G810gat,G811gat,G812gat,G813gat,G814gat,G815gat,G819gat,
G822gat,G825gat,G826gat,G827gat,G828gat,G829gat,G830gat,G831gat,G832gat,G833gat,
G834gat,G835gat,G836gat,G837gat,G838gat,G839gat,G840gat,G841gat,G842gat,G843gat,
G844gat,G845gat,G846gat,G847gat,G848gat,G849gat,G851gat,G852gat,G853gat,G854gat,
G855gat,G856gat,G857gat,G858gat,G859gat,G860gat,G861gat,G862gat,G867gat,G868gat,
G869gat,G870gat,G871gat,G872gat,G873gat,G875gat,G876gat,G877gat,muxed0,muxed1,
muxed2,muxed3,muxed4,muxed5,muxed6,muxed7,muxed8,muxed9,muxed10,muxed11,
muxed12,muxed13,muxed14,muxed15,muxed16,muxed17,muxed18,muxed19,muxed20,muxed21,
muxed22,muxed23,muxed24,muxed25,muxed26,muxed27,muxed28,muxed29,muxed30,muxed31,
muxed32,muxed33,muxed34,muxed35,muxed36,muxed37,muxed38,muxed39,muxed40,muxed41,
muxed42,muxed43,muxed44,muxed45,muxed46,muxed47,muxed48,muxed49,muxed50,muxed51,
muxed52,muxed53,muxed54,muxed55,muxed56,muxed57,muxed58,muxed59,muxed60,muxed61,
muxed62,muxed63,muxed64,muxed65,muxed66,muxed67,muxed68,muxed69,muxed70,muxed71,
muxed72,muxed73,muxed74,muxed75,muxed76,muxed77,muxed78,muxed79,muxed80,muxed81,
muxed82,muxed83,muxed84,muxed85,muxed86,muxed87,muxed88,muxed89,muxed90,muxed91,
muxed92,muxed93,muxed94,muxed95,muxed96,muxed97,muxed98,muxed99,muxed100,muxed101,
muxed102,muxed103,muxed104,muxed105,muxed106,muxed107,muxed108,muxed109,muxed110,muxed111,
muxed112,muxed113,muxed114,muxed115,muxed116,muxed117,muxed118,muxed119,muxed120,muxed121,
muxed122,muxed123,muxed124,muxed125,muxed126,muxed127,muxed128,muxed129,muxed130,muxed131,
muxed132,muxed133,muxed134,muxed135,muxed136,muxed137,muxed138,muxed139,muxed140,muxed141,
muxed142,muxed143,muxed144,muxed145,muxed146,muxed147,muxed148,muxed149,muxed150,muxed151,
muxed152,muxed153,muxed154,muxed155,muxed156,muxed157,muxed158,muxed159,muxed160,muxed161,
muxed162,muxed163,muxed164,muxed165,muxed166,muxed167,muxed168,muxed169,muxed170,muxed171,
muxed172,muxed173,muxed174,muxed175,muxed176,muxed177,muxed178,muxed179,muxed180,muxed181,
muxed182,muxed183,muxed184,muxed185,muxed186,muxed187,muxed188,muxed189,muxed190,muxed191,
muxed192,muxed193,muxed194,muxed195,muxed196,muxed197,muxed198,muxed199,muxed200,muxed201,
muxed202;
nand gate_0(G269gat,G1gat,G8gat,G13gat,muxed132);
nand gate_1(G270gat,G1gat,G26gat,G13gat,muxed132);
and gate_2(G273gat,G29gat,G36gat,G42gat);
and gate_3(G276gat,G1gat,G26gat,G51gat);
nand gate_4(G279gat,G1gat,G8gat,G51gat,muxed132);
nand gate_5(G280gat,G1gat,G8gat,G13gat,G55gat);
nand gate_6(G284gat,muxed43,G42gat,G68gat,G72gat);
nand gate_7(G285gat,G29gat,G68gat);
nand gate_8(G286gat,muxed43,G68gat,G74gat);
and gate_9(G287gat,G29gat,G75gat,G80gat);
and gate_10(G290gat,G29gat,G75gat,G42gat);
and gate_11(G291gat,G29gat,G36gat,G80gat);
and gate_12(G292gat,G29gat,G36gat,G42gat);
and gate_13(G293gat,muxed43,G75gat,G80gat);
and gate_14(G294gat,muxed43,G75gat,G42gat);
and gate_15(G295gat,muxed43,G36gat,G80gat);
and gate_16(G296gat,muxed43,G36gat,G42gat);
and gate_17(G297gat,G85gat,G86gat);
or gate_18(G298gat,G87gat,G88gat);
nand gate_19(G301gat,muxed81,G96gat);
or gate_20(G302gat,muxed81,G96gat);
nand gate_21(G303gat,G101gat,G106gat);
or gate_22(G304gat,G101gat,G106gat);
nand gate_23(G305gat,G111gat,G116gat);
or gate_24(G306gat,G111gat,G116gat);
nand gate_25(G307gat,G121gat,G126gat);
or gate_26(G308gat,G121gat,G126gat);
and gate_27(G309gat,G8gat,G138gat);
not gate_28(G310gat,G268gat);
and gate_29(G316gat,G51gat,G138gat);
and gate_30(G317gat,muxed132,G138gat);
and gate_31(G318gat,G152gat,G138gat);
nand gate_32(G319gat,muxed43,G156gat);
nor gate_33(G322gat,muxed132,G42gat);
and gate_34(G323gat,muxed132,G42gat);
nand gate_35(G324gat,G159gat,G165gat);
or gate_36(G325gat,G159gat,G165gat);
nand gate_37(G326gat,G171gat,G177gat);
or gate_38(G327gat,G171gat,G177gat);
nand gate_39(G328gat,G183gat,G189gat);
or gate_40(G329gat,G183gat,G189gat);
nand gate_41(G330gat,G195gat,G201gat);
or gate_42(G331gat,G195gat,G201gat);
and gate_43(G332gat,G210gat,muxed81);
and gate_44(G333gat,G210gat,G96gat);
and gate_45(G334gat,G210gat,G101gat);
and gate_46(G335gat,G210gat,G106gat);
and gate_47(G336gat,G210gat,G111gat);
and gate_48(G337gat,muxed69,G259gat);
and gate_49(G338gat,G210gat,G116gat);
and gate_50(G339gat,muxed69,G260gat);
and gate_51(G340gat,G210gat,G121gat);
and gate_52(G341gat,muxed69,G267gat);
not gate_53(G342gat,muxed108);
not gate_54(G343gat,G273gat);
or gate_55(G344gat,G270gat,G273gat);
not gate_56(G345gat,G276gat);
not gate_57(G346gat,G276gat);
not gate_58(G347gat,G279gat);
nor gate_59(G348gat,G280gat,G284gat);
or gate_60(G349gat,G280gat,G285gat);
or gate_61(G350gat,G280gat,G286gat);
not gate_62(G351gat,G293gat);
not gate_63(G352gat,G294gat);
not gate_64(G353gat,G295gat);
not gate_65(G354gat,G296gat);
nand gate_66(G355gat,G89gat,G298gat);
and gate_67(G356gat,G90gat,G298gat);
nand gate_68(G357gat,muxed91,G302gat);
nand gate_69(G360gat,G303gat,G304gat);
nand gate_70(G363gat,G305gat,G306gat);
nand gate_71(G366gat,G307gat,muxed173);
not gate_72(G369gat,G310gat);
nor gate_73(G375gat,G322gat,muxed159);
nand gate_74(G376gat,G324gat,G325gat);
nand gate_75(G379gat,G326gat,G327gat);
nand gate_76(G382gat,G328gat,muxed137);
nand gate_77(G385gat,G330gat,G331gat);
buf gate_78(G388gat,G290gat);
buf gate_79(G389gat,G291gat);
buf gate_80(G390gat,G292gat);
buf gate_81(G391gat,G297gat);
or gate_82(G392gat,G270gat,G343gat);
not gate_83(G393gat,G345gat);
not gate_84(G399gat,G346gat);
and gate_85(G400gat,G348gat,G73gat);
not gate_86(G401gat,G349gat);
not gate_87(G402gat,G350gat);
not gate_88(G403gat,G355gat);
not gate_89(G404gat,muxed90);
not gate_90(G405gat,muxed149);
and gate_91(G406gat,muxed90,muxed149);
not gate_92(G407gat,G363gat);
not gate_93(G408gat,G366gat);
and gate_94(G409gat,G363gat,G366gat);
nand gate_95(G410gat,G347gat,G352gat);
not gate_96(G411gat,G376gat);
not gate_97(G412gat,G379gat);
and gate_98(G413gat,G376gat,G379gat);
not gate_99(G414gat,G382gat);
not gate_100(G415gat,G385gat);
and gate_101(G416gat,G382gat,G385gat);
and gate_102(G417gat,G210gat,muxed27);
buf gate_103(G418gat,G342gat);
buf gate_104(G419gat,muxed92);
buf gate_105(G420gat,G351gat);
buf gate_106(G421gat,G353gat);
buf gate_107(G422gat,G354gat);
buf gate_108(G423gat,G356gat);
not gate_109(G424gat,G400gat);
and gate_110(G425gat,muxed171,G405gat);
and gate_111(G426gat,G407gat,G408gat);
and gate_112(G427gat,muxed55,G393gat,G55gat);
and gate_113(G432gat,G393gat,muxed132,G287gat);
nand gate_114(G437gat,G393gat,G287gat,G55gat);
nand gate_115(G442gat,muxed180,muxed43,G156gat,G393gat);
nand gate_116(G443gat,G393gat,muxed55,muxed132);
and gate_117(G444gat,G411gat,G412gat);
and gate_118(G445gat,G414gat,muxed9);
buf gate_119(G446gat,G392gat);
buf gate_120(G447gat,G399gat);
buf gate_121(G448gat,G401gat);
buf gate_122(G449gat,G402gat);
buf gate_123(G450gat,G403gat);
not gate_124(G451gat,G424gat);
nor gate_125(G460gat,muxed88,muxed18);
nor gate_126(G463gat,muxed147,G426gat);
nand gate_127(G466gat,muxed188,G410gat);
and gate_128(G475gat,G143gat,G427gat);
and gate_129(G476gat,G310gat,G432gat);
and gate_130(G477gat,G146gat,G427gat);
and gate_131(G478gat,G310gat,G432gat);
and gate_132(G479gat,G149gat,G427gat);
and gate_133(G480gat,G310gat,G432gat);
and gate_134(G481gat,G153gat,G427gat);
and gate_135(G482gat,G310gat,G432gat);
nand gate_136(G483gat,muxed64,G1gat);
or gate_137(G488gat,muxed27,G437gat);
or gate_138(G489gat,muxed27,G437gat);
or gate_139(G490gat,muxed27,G437gat);
or gate_140(G491gat,muxed27,G437gat);
nor gate_141(G492gat,G413gat,G444gat);
nor gate_142(G495gat,G416gat,G445gat);
nand gate_143(G498gat,G130gat,muxed87);
or gate_144(G499gat,G130gat,muxed87);
nand gate_145(G500gat,G463gat,G135gat);
or gate_146(G501gat,G463gat,G135gat);
and gate_147(G502gat,muxed81,G466gat);
nor gate_148(G503gat,G475gat,G476gat);
and gate_149(G504gat,G96gat,G466gat);
nor gate_150(G505gat,G477gat,G478gat);
and gate_151(G506gat,G101gat,G466gat);
nor gate_152(G507gat,G479gat,G480gat);
and gate_153(G508gat,G106gat,G466gat);
nor gate_154(G509gat,G481gat,G482gat);
and gate_155(G510gat,G143gat,muxed193);
and gate_156(G511gat,G111gat,G466gat);
and gate_157(G512gat,G146gat,muxed193);
and gate_158(G513gat,G116gat,G466gat);
and gate_159(G514gat,G149gat,muxed193);
and gate_160(G515gat,G121gat,G466gat);
and gate_161(G516gat,G153gat,muxed193);
and gate_162(G517gat,G126gat,G466gat);
nand gate_163(G518gat,G130gat,G492gat);
or gate_164(G519gat,G130gat,G492gat);
nand gate_165(G520gat,G495gat,G207gat);
or gate_166(G521gat,G495gat,G207gat);
and gate_167(G522gat,G451gat,G159gat);
and gate_168(G523gat,G451gat,G165gat);
and gate_169(G524gat,G451gat,G171gat);
and gate_170(G525gat,G451gat,G177gat);
and gate_171(G526gat,G451gat,G183gat);
nand gate_172(G527gat,G451gat,G189gat);
nand gate_173(G528gat,G451gat,G195gat);
nand gate_174(G529gat,G451gat,G201gat);
nand gate_175(G530gat,G498gat,muxed85);
nand gate_176(G533gat,G500gat,G501gat);
nor gate_177(G536gat,G309gat,muxed166);
nor gate_178(G537gat,muxed140,G504gat);
nor gate_179(G538gat,G317gat,G506gat);
nor gate_180(G539gat,G318gat,G508gat);
nor gate_181(G540gat,G510gat,G511gat);
nor gate_182(G541gat,G512gat,G513gat);
nor gate_183(G542gat,G514gat,G515gat);
nor gate_184(G543gat,muxed127,G517gat);
nand gate_185(G544gat,muxed182,G519gat);
nand gate_186(G547gat,muxed89,G521gat);
not gate_187(G550gat,muxed46);
not gate_188(G551gat,muxed56);
and gate_189(G552gat,muxed46,muxed56);
nand gate_190(G553gat,G536gat,muxed35);
nand gate_191(G557gat,muxed152,G505gat);
nand gate_192(G561gat,muxed58,muxed178);
nand gate_193(G565gat,muxed175,muxed72);
nand gate_194(G569gat,G488gat,G540gat);
nand gate_195(G573gat,G489gat,G541gat);
nand gate_196(G577gat,muxed141,muxed83);
nand gate_197(G581gat,muxed176,muxed48);
not gate_198(G585gat,muxed164);
not gate_199(G586gat,G547gat);
and gate_200(G587gat,muxed164,G547gat);
and gate_201(G588gat,G550gat,muxed67);
and gate_202(G589gat,G585gat,G586gat);
nand gate_203(G590gat,G553gat,G159gat);
or gate_204(G593gat,G553gat,G159gat);
and gate_205(G596gat,muxed93,G553gat);
nand gate_206(G597gat,muxed155,G165gat);
or gate_207(G600gat,muxed155,G165gat);
and gate_208(G605gat,muxed93,muxed155);
nand gate_209(G606gat,muxed57,G171gat);
or gate_210(G609gat,muxed57,G171gat);
and gate_211(G615gat,muxed93,muxed57);
nand gate_212(G616gat,muxed174,G177gat);
or gate_213(G619gat,muxed174,G177gat);
and gate_214(G624gat,muxed93,muxed174);
nand gate_215(G625gat,G569gat,G183gat);
or gate_216(G628gat,G569gat,G183gat);
and gate_217(G631gat,muxed93,G569gat);
nand gate_218(G632gat,muxed95,G189gat);
or gate_219(G635gat,muxed95,G189gat);
and gate_220(G640gat,muxed93,muxed95);
nand gate_221(G641gat,muxed40,G195gat);
or gate_222(G644gat,muxed40,G195gat);
and gate_223(G650gat,muxed93,muxed40);
nand gate_224(G651gat,muxed194,G201gat);
or gate_225(G654gat,muxed194,G201gat);
and gate_226(G659gat,muxed93,muxed194);
nor gate_227(G660gat,G552gat,muxed66);
nor gate_228(G661gat,G587gat,G589gat);
not gate_229(G662gat,G590gat);
and gate_230(G665gat,G593gat,G590gat);
nor gate_231(G669gat,G596gat,G522gat);
not gate_232(G670gat,muxed138);
and gate_233(G673gat,muxed167,muxed138);
nor gate_234(G677gat,muxed73,G523gat);
not gate_235(G678gat,G606gat);
and gate_236(G682gat,G609gat,G606gat);
nor gate_237(G686gat,G615gat,G524gat);
not gate_238(G687gat,G616gat);
and gate_239(G692gat,G619gat,G616gat);
nor gate_240(G696gat,muxed172,G525gat);
not gate_241(G697gat,G625gat);
and gate_242(G700gat,G628gat,G625gat);
nor gate_243(G704gat,G631gat,G526gat);
not gate_244(G705gat,G632gat);
and gate_245(G708gat,muxed0,G632gat);
nor gate_246(G712gat,G337gat,muxed94);
not gate_247(G713gat,G641gat);
and gate_248(G717gat,G644gat,G641gat);
nor gate_249(G721gat,muxed79,muxed38);
not gate_250(G722gat,muxed129);
and gate_251(G727gat,G654gat,muxed129);
nor gate_252(G731gat,G341gat,muxed45);
nand gate_253(G732gat,G654gat,G261gat);
nand gate_254(G733gat,G644gat,G654gat,G261gat);
nand gate_255(G734gat,muxed0,G644gat,G654gat,G261gat);
not gate_256(G735gat,muxed202);
and gate_257(G736gat,G228gat,G665gat);
and gate_258(G737gat,G237gat,muxed202);
not gate_259(G738gat,G670gat);
and gate_260(G739gat,G228gat,muxed135);
and gate_261(G740gat,G237gat,G670gat);
not gate_262(G741gat,G678gat);
and gate_263(G742gat,G228gat,G682gat);
and gate_264(G743gat,G237gat,G678gat);
not gate_265(G744gat,G687gat);
and gate_266(G745gat,G228gat,muxed42);
and gate_267(G746gat,G237gat,G687gat);
not gate_268(G747gat,G697gat);
and gate_269(G748gat,G228gat,G700gat);
and gate_270(G749gat,G237gat,G697gat);
not gate_271(G750gat,G705gat);
and gate_272(G751gat,G228gat,muxed191);
and gate_273(G752gat,G237gat,G705gat);
not gate_274(G753gat,muxed153);
and gate_275(G754gat,G228gat,G717gat);
and gate_276(G755gat,G237gat,muxed153);
not gate_277(G756gat,G722gat);
nor gate_278(G757gat,muxed154,G261gat);
and gate_279(G758gat,muxed154,G261gat);
and gate_280(G759gat,G228gat,muxed154);
and gate_281(G760gat,G237gat,G722gat);
nand gate_282(G761gat,G644gat,G722gat);
nand gate_283(G762gat,muxed0,muxed153);
nand gate_284(G763gat,muxed0,G644gat,G722gat);
nand gate_285(G764gat,G609gat,G687gat);
nand gate_286(G765gat,muxed167,G678gat);
nand gate_287(G766gat,muxed167,G609gat,G687gat);
buf gate_288(G767gat,G660gat);
buf gate_289(G768gat,G661gat);
nor gate_290(G769gat,G736gat,G737gat);
nor gate_291(G770gat,G739gat,G740gat);
nor gate_292(G771gat,G742gat,G743gat);
nor gate_293(G772gat,G745gat,G746gat);
nand gate_294(G773gat,muxed151,muxed11,G763gat,G734gat);
nor gate_295(G777gat,G748gat,G749gat);
nand gate_296(G778gat,G753gat,G761gat,G733gat);
nor gate_297(G781gat,G751gat,muxed199);
nand gate_298(G782gat,G756gat,G732gat);
nor gate_299(G785gat,G754gat,muxed197);
nor gate_300(G786gat,muxed165,G758gat);
nor gate_301(G787gat,muxed126,G760gat);
nor gate_302(G788gat,G700gat,muxed10);
and gate_303(G789gat,G700gat,muxed10);
nor gate_304(G790gat,muxed191,G778gat);
and gate_305(G791gat,muxed191,G778gat);
nor gate_306(G792gat,G717gat,muxed54);
and gate_307(G793gat,G717gat,muxed54);
and gate_308(G794gat,G219gat,muxed184);
nand gate_309(G795gat,G628gat,muxed10);
nand gate_310(G796gat,muxed8,G747gat);
nor gate_311(G802gat,G788gat,G789gat);
nor gate_312(G803gat,muxed201,G791gat);
nor gate_313(G804gat,G792gat,G793gat);
nor gate_314(G805gat,muxed22,muxed160);
nor gate_315(G806gat,muxed42,muxed7);
and gate_316(G807gat,muxed42,muxed7);
and gate_317(G808gat,G219gat,G802gat);
and gate_318(G809gat,G219gat,muxed200);
and gate_319(G810gat,G219gat,G804gat);
nand gate_320(G811gat,G805gat,muxed124,muxed44,G529gat);
nand gate_321(G812gat,G619gat,muxed7);
nand gate_322(G813gat,G609gat,G619gat,muxed7);
nand gate_323(G814gat,muxed167,G609gat,G619gat,muxed7);
nand gate_324(G815gat,G738gat,G765gat,G766gat,muxed5);
nand gate_325(G819gat,G741gat,G764gat,G813gat);
nand gate_326(G822gat,G744gat,G812gat);
nor gate_327(G825gat,G806gat,G807gat);
nor gate_328(G826gat,muxed29,G808gat);
nor gate_329(G827gat,G336gat,G809gat);
nor gate_330(G828gat,G338gat,G810gat);
not gate_331(G829gat,muxed122);
nor gate_332(G830gat,G665gat,muxed97);
and gate_333(G831gat,G665gat,muxed97);
nor gate_334(G832gat,muxed135,G819gat);
and gate_335(G833gat,muxed135,G819gat);
nor gate_336(G834gat,G682gat,muxed12);
and gate_337(G835gat,G682gat,muxed12);
and gate_338(G836gat,G219gat,G825gat);
nand gate_339(G837gat,G826gat,G777gat,muxed20);
nand gate_340(G838gat,G827gat,G781gat,G712gat,G527gat);
nand gate_341(G839gat,G828gat,G785gat,muxed80,G528gat);
not gate_342(G840gat,muxed130);
nand gate_343(G841gat,muxed97,G593gat);
nor gate_344(G842gat,G830gat,G831gat);
nor gate_345(G843gat,G832gat,muxed23);
nor gate_346(G844gat,muxed16,G835gat);
nor gate_347(G845gat,G334gat,muxed101);
not gate_348(G846gat,G837gat);
not gate_349(G847gat,G838gat);
not gate_350(G848gat,muxed34);
and gate_351(G849gat,G735gat,muxed2);
buf gate_352(G850gat,muxed143);
and gate_353(G851gat,G219gat,G842gat);
and gate_354(G852gat,G219gat,muxed21);
and gate_355(G853gat,G219gat,G844gat);
nand gate_356(G854gat,muxed99,G772gat,muxed170);
not gate_357(G855gat,G846gat);
not gate_358(G856gat,G847gat);
not gate_359(G857gat,muxed32);
not gate_360(G858gat,muxed1);
nor gate_361(G859gat,muxed186,G851gat);
nor gate_362(G860gat,G332gat,muxed19);
nor gate_363(G861gat,G333gat,G853gat);
not gate_364(G862gat,muxed98);
buf gate_365(G863gat,muxed157);
buf gate_366(G864gat,G856gat);
buf gate_367(G865gat,muxed30);
buf gate_368(G866gat,G858gat);
nand gate_369(G867gat,G859gat,G769gat,G669gat);
nand gate_370(G868gat,muxed119,G770gat,muxed198);
nand gate_371(G869gat,G861gat,G771gat,G686gat);
not gate_372(G870gat,G862gat);
not gate_373(G871gat,G867gat);
not gate_374(G872gat,muxed15);
not gate_375(G873gat,G869gat);
buf gate_376(G874gat,G870gat);
not gate_377(G875gat,G871gat);
not gate_378(G876gat,muxed76);
not gate_379(G877gat,G873gat);
buf gate_380(G878gat,G875gat);
buf gate_381(G879gat,G876gat);
buf gate_382(G880gat,G877gat);
assign muxed0 = keyinput0 ? muxed24 : muxed1;
assign muxed1 = keyinput1 ? muxed102 : G678gat;
assign muxed2 = keyinput2 ? muxed96 : muxed147;
assign muxed3 = keyinput3 ? G573gat : muxed96;
assign muxed4 = keyinput4 ? G815gat : muxed98;
assign muxed5 = keyinput5 ? muxed179 : muxed0;
assign muxed6 = keyinput6 ? G539gat : muxed179;
assign muxed7 = keyinput7 ? muxed31 : G346gat;
assign muxed8 = keyinput8 ? G795gat : muxed200;
assign muxed9 = keyinput9 ? G415gat : G795gat;
assign muxed10 = keyinput10 ? G773gat : G353gat;
assign muxed11 = keyinput11 ? G762gat : G403gat;
assign muxed12 = keyinput12 ? G822gat : G762gat;
assign muxed13 = keyinput13 ? muxed150 : muxed76;
assign muxed14 = keyinput14 ? G872gat : muxed83;
assign muxed15 = keyinput15 ? muxed70 : muxed44;
assign muxed16 = keyinput16 ? G834gat : muxed70;
assign muxed17 = keyinput17 ? G860gat : muxed130;
assign muxed18 = keyinput18 ? G425gat : G860gat;
assign muxed19 = keyinput19 ? G852gat : G873gat;
assign muxed20 = keyinput20 ? G704gat : G852gat;
assign muxed21 = keyinput21 ? G843gat : G644gat;
assign muxed22 = keyinput22 ? muxed190 : G843gat;
assign muxed23 = keyinput23 ? muxed134 : G819gat;
assign muxed24 = keyinput24 ? G635gat : muxed134;
assign muxed25 = keyinput25 ? muxed136 : G334gat;
assign muxed26 = keyinput26 ? muxed86 : muxed143;
assign muxed27 = keyinput27 ? G369gat : muxed28;
assign muxed28 = keyinput28 ? G865gat : muxed40;
assign muxed29 = keyinput29 ? G335gat : G865gat;
assign muxed30 = keyinput30 ? G857gat : G749gat;
assign muxed31 = keyinput31 ? G796gat : G857gat;
assign muxed32 = keyinput32 ? G848gat : G812gat;
assign muxed33 = keyinput33 ? muxed177 : G848gat;
assign muxed34 = keyinput34 ? G839gat : G764gat;
assign muxed35 = keyinput35 ? muxed100 : G839gat;
assign muxed36 = keyinput36 ? muxed78 : G766gat;
assign muxed37 = keyinput37 ? G542gat : muxed78;
assign muxed38 = keyinput38 ? muxed103 : G505gat;
assign muxed39 = keyinput39 ? muxed68 : muxed103;
assign muxed40 = keyinput40 ? G577gat : muxed182;
assign muxed41 = keyinput41 ? G490gat : G348gat;
assign muxed42 = keyinput42 ? G692gat : G490gat;
assign muxed43 = keyinput43 ? G59gat : muxed44;
assign muxed44 = keyinput44 ? G731gat : G303gat;
assign muxed45 = keyinput45 ? G659gat : G451gat;
assign muxed46 = keyinput46 ? muxed84 : G659gat;
assign muxed47 = keyinput47 ? G581gat : G819gat;
assign muxed48 = keyinput48 ? G543gat : G481gat;
assign muxed49 = keyinput49 ? muxed142 : G543gat;
assign muxed50 = keyinput50 ? muxed106 : G741gat;
assign muxed51 = keyinput51 ? G538gat : muxed106;
assign muxed52 = keyinput52 ? muxed120 : muxed188;
assign muxed53 = keyinput53 ? muxed131 : muxed66;
assign muxed54 = keyinput54 ? G782gat : muxed131;
assign muxed55 = keyinput55 ? G319gat : G577gat;
assign muxed56 = keyinput56 ? G533gat : muxed57;
assign muxed57 = keyinput57 ? muxed59 : G317gat;
assign muxed58 = keyinput58 ? muxed133 : G705gat;
assign muxed59 = keyinput59 ? muxed65 : muxed133;
assign muxed60 = keyinput60 ? muxed107 : G304gat;
assign muxed61 = keyinput61 ? muxed110 : G333gat;
assign muxed62 = keyinput62 ? G483gat : G661gat;
assign muxed63 = keyinput63 ? G503gat : G483gat;
assign muxed64 = keyinput64 ? muxed53 : muxed38;
assign muxed65 = keyinput65 ? G561gat : muxed53;
assign muxed66 = keyinput66 ? G588gat : G573gat;
assign muxed67 = keyinput67 ? G551gat : muxed29;
assign muxed68 = keyinput68 ? G836gat : G551gat;
assign muxed69 = keyinput69 ? G255gat : muxed70;
assign muxed70 = keyinput70 ? muxed195 : muxed57;
assign muxed71 = keyinput71 ? G677gat : muxed200;
assign muxed72 = keyinput72 ? G509gat : G677gat;
assign muxed73 = keyinput73 ? muxed144 : G332gat;
assign muxed74 = keyinput74 ? muxed41 : muxed144;
assign muxed75 = keyinput75 ? muxed148 : G585gat;
assign muxed76 = keyinput76 ? muxed82 : G332gat;
assign muxed77 = keyinput77 ? muxed37 : muxed84;
assign muxed78 = keyinput78 ? G721gat : G432gat;
assign muxed79 = keyinput79 ? G339gat : muxed0;
assign muxed80 = keyinput80 ? muxed36 : G339gat;
assign muxed81 = keyinput81 ? G91gat : muxed82;
assign muxed82 = keyinput82 ? muxed14 : G749gat;
assign muxed83 = keyinput83 ? muxed77 : G704gat;
assign muxed84 = keyinput84 ? G530gat : G552gat;
assign muxed85 = keyinput85 ? G499gat : G735gat;
assign muxed86 = keyinput86 ? G597gat : G499gat;
assign muxed87 = keyinput87 ? G460gat : G526gat;
assign muxed88 = keyinput88 ? G406gat : G479gat;
assign muxed89 = keyinput89 ? G520gat : G406gat;
assign muxed90 = keyinput90 ? G357gat : G533gat;
assign muxed91 = keyinput91 ? G301gat : G772gat;
assign muxed92 = keyinput92 ? G344gat : G301gat;
assign muxed93 = keyinput93 ? G246gat : muxed94;
assign muxed94 = keyinput94 ? G640gat : muxed73;
assign muxed95 = keyinput95 ? muxed3 : G867gat;
assign muxed96 = keyinput96 ? G841gat : G819gat;
assign muxed97 = keyinput97 ? muxed4 : muxed191;
assign muxed98 = keyinput98 ? muxed169 : G415gat;
assign muxed99 = keyinput99 ? G845gat : G872gat;
assign muxed100 = keyinput100 ? muxed63 : G845gat;
assign muxed101 = keyinput101 ? muxed39 : G788gat;
assign muxed102 = keyinput102 ? G849gat : muxed39;
assign muxed103 = keyinput103 ? muxed116 : G273gat;
assign muxed104 = keyinput104 ? G17gat : muxed133;
assign muxed105 = keyinput105 ? muxed51 : muxed134;
assign muxed106 = keyinput106 ? muxed60 : G348gat;
assign muxed107 = keyinput107 ? muxed192 : G319gat;
assign muxed108 = keyinput108 ? G269gat : muxed192;
assign muxed109 = keyinput109 ? muxed61 : muxed194;
assign muxed110 = keyinput110 ? muxed187 : muxed103;
assign muxed111 = keyinput111 ? G417gat : muxed187;
assign muxed112 = keyinput112 ? muxed189 : G843gat;
assign muxed113 = keyinput113 ? muxed158 : G809gat;
assign muxed114 = keyinput114 ? muxed168 : muxed158;
assign muxed115 = keyinput115 ? G323gat : muxed160;
assign muxed116 = keyinput116 ? G650gat : G323gat;
assign muxed117 = keyinput117 ? muxed47 : muxed195;
assign muxed118 = keyinput118 ? muxed196 : G508gat;
assign muxed119 = keyinput119 ? muxed17 : muxed199;
assign muxed120 = keyinput120 ? muxed123 : muxed17;
assign muxed121 = keyinput121 ? G829gat : muxed182;
assign muxed122 = keyinput122 ? G811gat : G525gat;
assign muxed123 = keyinput123 ? muxed62 : G811gat;
assign muxed124 = keyinput124 ? G787gat : G842gat;
assign muxed125 = keyinput125 ? muxed161 : G787gat;
assign muxed126 = keyinput126 ? G759gat : G347gat;
assign muxed127 = keyinput127 ? muxed50 : G759gat;
assign muxed128 = keyinput128 ? G727gat : muxed202;
assign muxed129 = keyinput129 ? G651gat : muxed137;
assign muxed130 = keyinput130 ? muxed181 : muxed131;
assign muxed131 = keyinput131 ? G443gat : muxed21;
assign muxed132 = keyinput132 ? muxed104 : G789gat;
assign muxed133 = keyinput133 ? muxed105 : G717gat;
assign muxed134 = keyinput134 ? G833gat : G412gat;
assign muxed135 = keyinput135 ? muxed25 : muxed15;
assign muxed136 = keyinput136 ? G673gat : G296gat;
assign muxed137 = keyinput137 ? G329gat : G673gat;
assign muxed138 = keyinput138 ? muxed26 : muxed35;
assign muxed139 = keyinput139 ? G840gat : G593gat;
assign muxed140 = keyinput140 ? G316gat : muxed141;
assign muxed141 = keyinput141 ? muxed49 : G400gat;
assign muxed142 = keyinput142 ? muxed74 : G529gat;
assign muxed143 = keyinput143 ? muxed139 : muxed74;
assign muxed144 = keyinput144 ? G605gat : G293gat;
assign muxed145 = keyinput145 ? muxed156 : muxed0;
assign muxed146 = keyinput146 ? muxed75 : muxed169;
assign muxed147 = keyinput147 ? G409gat : muxed75;
assign muxed148 = keyinput148 ? muxed13 : muxed28;
assign muxed149 = keyinput149 ? G360gat : muxed13;
assign muxed150 = keyinput150 ? G557gat : muxed12;
assign muxed151 = keyinput151 ? G750gat : G557gat;
assign muxed152 = keyinput152 ? G537gat : muxed73;
assign muxed153 = keyinput153 ? G713gat : G537gat;
assign muxed154 = keyinput154 ? muxed185 : muxed155;
assign muxed155 = keyinput155 ? muxed145 : G405gat;
assign muxed156 = keyinput156 ? muxed114 : muxed123;
assign muxed157 = keyinput157 ? G855gat : muxed114;
assign muxed158 = keyinput158 ? G375gat : muxed159;
assign muxed159 = keyinput159 ? muxed115 : G280gat;
assign muxed160 = keyinput160 ? muxed125 : muxed62;
assign muxed161 = keyinput161 ? muxed183 : muxed99;
assign muxed162 = keyinput162 ? G518gat : muxed183;
assign muxed163 = keyinput163 ? G786gat : muxed186;
assign muxed164 = keyinput164 ? G544gat : G786gat;
assign muxed165 = keyinput165 ? G757gat : G759gat;
assign muxed166 = keyinput166 ? G502gat : G757gat;
assign muxed167 = keyinput167 ? G600gat : muxed168;
assign muxed168 = keyinput168 ? muxed146 : muxed78;
assign muxed169 = keyinput169 ? G854gat : G828gat;
assign muxed170 = keyinput170 ? G696gat : muxed101;
assign muxed171 = keyinput171 ? G404gat : G696gat;
assign muxed172 = keyinput172 ? G624gat : muxed142;
assign muxed173 = keyinput173 ? G308gat : G624gat;
assign muxed174 = keyinput174 ? G565gat : muxed125;
assign muxed175 = keyinput175 ? muxed33 : G513gat;
assign muxed176 = keyinput176 ? G491gat : muxed33;
assign muxed177 = keyinput177 ? muxed6 : G635gat;
assign muxed178 = keyinput178 ? G507gat : muxed6;
assign muxed179 = keyinput179 ? G814gat : G539gat;
assign muxed180 = keyinput180 ? muxed113 : muxed181;
assign muxed181 = keyinput181 ? muxed121 : G269gat;
assign muxed182 = keyinput182 ? muxed162 : muxed92;
assign muxed183 = keyinput183 ? G794gat : muxed75;
assign muxed184 = keyinput184 ? muxed163 : G659gat;
assign muxed185 = keyinput185 ? muxed128 : muxed163;
assign muxed186 = keyinput186 ? muxed111 : G505gat;
assign muxed187 = keyinput187 ? muxed52 : G813gat;
assign muxed188 = keyinput188 ? muxed112 : muxed173;
assign muxed189 = keyinput189 ? G442gat : muxed7;
assign muxed190 = keyinput190 ? G340gat : G442gat;
assign muxed191 = keyinput191 ? G708gat : muxed192;
assign muxed192 = keyinput192 ? G516gat : G331gat;
assign muxed193 = keyinput193 ? muxed109 : G644gat;
assign muxed194 = keyinput194 ? muxed117 : G677gat;
assign muxed195 = keyinput195 ? muxed118 : muxed17;
assign muxed196 = keyinput196 ? G868gat : muxed153;
assign muxed197 = keyinput197 ? G755gat : G868gat;
assign muxed198 = keyinput198 ? muxed71 : G326gat;
assign muxed199 = keyinput199 ? G752gat : muxed71;
assign muxed200 = keyinput200 ? G803gat : muxed160;
assign muxed201 = keyinput201 ? G790gat : muxed175;
assign muxed202 = keyinput202 ? G662gat : G790gat;
endmodule
