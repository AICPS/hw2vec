// Verilog File 
module top (G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,
G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,
G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,
G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat,G223gat,G329gat,G370gat,
G421gat,G430gat,G431gat,G432gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,
keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,
keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,
keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,keyinput35,
keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,keyinput45,
keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,keyinput55,
keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,keyinput65,
keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,keyinput75,
keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,keyinput85,
keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,keyinput95,
keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101);

input G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,
G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,
G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,
G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat,keyinput0,keyinput1,keyinput2,
keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,
keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,
keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,
keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,
keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,
keyinput53,keyinput54,keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,
keyinput63,keyinput64,keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,
keyinput73,keyinput74,keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,
keyinput83,keyinput84,keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,
keyinput93,keyinput94,keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101;

output G223gat,G329gat,G370gat,G421gat,G430gat,G431gat,G432gat;

wire G118gat,G119gat,G122gat,G123gat,G126gat,G127gat,G130gat,G131gat,G134gat,
G135gat,G138gat,G139gat,G142gat,G143gat,G146gat,G147gat,G150gat,G151gat,G154gat,
G157gat,G158gat,G159gat,G162gat,G165gat,G168gat,G171gat,G174gat,G177gat,G180gat,
G183gat,G184gat,G185gat,G186gat,G187gat,G188gat,G189gat,G190gat,G191gat,G192gat,
G193gat,G194gat,G195gat,G196gat,G197gat,G198gat,G199gat,G203gat,G213gat,G224gat,
G227gat,G230gat,G233gat,G236gat,G239gat,G242gat,G243gat,G246gat,G247gat,G250gat,
G251gat,G254gat,G255gat,G256gat,G257gat,G258gat,G259gat,G260gat,G263gat,G264gat,
G267gat,G270gat,G273gat,G276gat,G279gat,G282gat,G285gat,G288gat,G289gat,G290gat,
G291gat,G292gat,G293gat,G294gat,G295gat,G296gat,G300gat,G301gat,G302gat,G303gat,
G304gat,G305gat,G306gat,G307gat,G308gat,G309gat,G319gat,G330gat,G331gat,G332gat,
G333gat,G334gat,G335gat,G336gat,G337gat,G338gat,G339gat,G340gat,G341gat,G342gat,
G343gat,G344gat,G345gat,G346gat,G347gat,G348gat,G349gat,G350gat,G351gat,G352gat,
G353gat,G354gat,G355gat,G356gat,G357gat,G360gat,G371gat,G372gat,G373gat,G374gat,
G375gat,G376gat,G377gat,G378gat,G379gat,G380gat,G381gat,G386gat,G393gat,G399gat,
G404gat,G407gat,G411gat,G414gat,G415gat,G416gat,G417gat,G418gat,G419gat,G420gat,
G422gat,G425gat,G428gat,G429gat,muxed0,muxed1,muxed2,muxed3,muxed4,muxed5,
muxed6,muxed7,muxed8,muxed9,muxed10,muxed11,muxed12,muxed13,muxed14,muxed15,
muxed16,muxed17,muxed18,muxed19,muxed20,muxed21,muxed22,muxed23,muxed24,muxed25,
muxed26,muxed27,muxed28,muxed29,muxed30,muxed31,muxed32,muxed33,muxed34,muxed35,
muxed36,muxed37,muxed38,muxed39,muxed40,muxed41,muxed42,muxed43,muxed44,muxed45,
muxed46,muxed47,muxed48,muxed49,muxed50,muxed51,muxed52,muxed53,muxed54,muxed55,
muxed56,muxed57,muxed58,muxed59,muxed60,muxed61,muxed62,muxed63,muxed64,muxed65,
muxed66,muxed67,muxed68,muxed69,muxed70,muxed71,muxed72,muxed73,muxed74,muxed75,
muxed76,muxed77,muxed78,muxed79,muxed80,muxed81,muxed82,muxed83,muxed84,muxed85,
muxed86,muxed87,muxed88,muxed89,muxed90,muxed91,muxed92,muxed93,muxed94,muxed95,
muxed96,muxed97,muxed98,muxed99,muxed100,muxed101;
not gate_0(G118gat,G1gat);
not gate_1(G119gat,G4gat);
not gate_2(G122gat,G11gat);
not gate_3(G123gat,muxed76);
not gate_4(G126gat,G24gat);
not gate_5(G127gat,G30gat);
not gate_6(G130gat,G37gat);
not gate_7(G131gat,G43gat);
not gate_8(G134gat,G50gat);
not gate_9(G135gat,G56gat);
not gate_10(G138gat,G63gat);
not gate_11(G139gat,G69gat);
not gate_12(G142gat,G76gat);
not gate_13(G143gat,G82gat);
not gate_14(G146gat,G89gat);
not gate_15(G147gat,G95gat);
not gate_16(G150gat,G102gat);
not gate_17(G151gat,G108gat);
nand gate_18(G154gat,G118gat,G4gat);
nor gate_19(G157gat,G8gat,G119gat);
nor gate_20(G158gat,G14gat,G119gat);
nand gate_21(G159gat,G122gat,muxed76);
nand gate_22(G162gat,G126gat,G30gat);
nand gate_23(G165gat,muxed79,G43gat);
nand gate_24(G168gat,muxed87,G56gat);
nand gate_25(G171gat,G138gat,G69gat);
nand gate_26(G174gat,muxed92,G82gat);
nand gate_27(G177gat,G146gat,G95gat);
nand gate_28(G180gat,G150gat,G108gat);
nor gate_29(G183gat,G21gat,muxed88);
nor gate_30(G184gat,G27gat,muxed88);
nor gate_31(G185gat,G34gat,G127gat);
nor gate_32(G186gat,G40gat,G127gat);
nor gate_33(G187gat,G47gat,G131gat);
nor gate_34(G188gat,G53gat,G131gat);
nor gate_35(G189gat,G60gat,G135gat);
nor gate_36(G190gat,G66gat,G135gat);
nor gate_37(G191gat,muxed26,G139gat);
nor gate_38(G192gat,G79gat,G139gat);
nor gate_39(G193gat,G86gat,G143gat);
nor gate_40(G194gat,G92gat,G143gat);
nor gate_41(G195gat,G99gat,G147gat);
nor gate_42(G196gat,G105gat,G147gat);
nor gate_43(G197gat,G112gat,G151gat);
nor gate_44(G198gat,G115gat,G151gat);
and gate_45(G199gat,G154gat,muxed72,G162gat,G165gat,G168gat,muxed46,muxed49,G177gat,muxed43);
not gate_46(G203gat,G199gat);
not gate_47(G213gat,G199gat);
not gate_48(G223gat,G199gat);
xor gate_49(G224gat,G203gat,G154gat);
xor gate_50(G227gat,G203gat,muxed72);
xor gate_51(G230gat,G203gat,G162gat);
xor gate_52(G233gat,G203gat,G165gat);
xor gate_53(G236gat,G203gat,G168gat);
xor gate_54(G239gat,G203gat,muxed46);
nand gate_55(G242gat,G1gat,G213gat);
xor gate_56(G243gat,G203gat,muxed49);
nand gate_57(G246gat,G213gat,G11gat);
xor gate_58(G247gat,G203gat,G177gat);
nand gate_59(G250gat,G213gat,G24gat);
xor gate_60(G251gat,G203gat,muxed43);
nand gate_61(G254gat,G213gat,G37gat);
nand gate_62(G255gat,G213gat,G50gat);
nand gate_63(G256gat,G213gat,G63gat);
nand gate_64(G257gat,G213gat,G76gat);
nand gate_65(G258gat,G213gat,G89gat);
nand gate_66(G259gat,G213gat,G102gat);
nand gate_67(G260gat,G224gat,G157gat);
nand gate_68(G263gat,G224gat,G158gat);
nand gate_69(G264gat,muxed71,G183gat);
nand gate_70(G267gat,G230gat,G185gat);
nand gate_71(G270gat,muxed21,G187gat);
nand gate_72(G273gat,muxed90,G189gat);
nand gate_73(G276gat,G239gat,muxed38);
nand gate_74(G279gat,muxed48,G193gat);
nand gate_75(G282gat,G247gat,muxed29);
nand gate_76(G285gat,G251gat,G197gat);
nand gate_77(G288gat,muxed71,muxed86);
nand gate_78(G289gat,G230gat,G186gat);
nand gate_79(G290gat,muxed21,muxed19);
nand gate_80(G291gat,muxed90,G190gat);
nand gate_81(G292gat,G239gat,muxed84);
nand gate_82(G293gat,muxed48,G194gat);
nand gate_83(G294gat,G247gat,G196gat);
nand gate_84(G295gat,G251gat,G198gat);
and gate_85(G296gat,G260gat,G264gat,muxed37,G270gat,muxed62,G276gat,G279gat,G282gat,G285gat);
not gate_86(G300gat,G263gat);
not gate_87(G301gat,muxed67);
not gate_88(G302gat,G289gat);
not gate_89(G303gat,muxed45);
not gate_90(G304gat,G291gat);
not gate_91(G305gat,G292gat);
not gate_92(G306gat,muxed47);
not gate_93(G307gat,muxed68);
not gate_94(G308gat,G295gat);
not gate_95(G309gat,G296gat);
not gate_96(G319gat,G296gat);
not gate_97(G329gat,G296gat);
xor gate_98(G330gat,muxed95,G260gat);
xor gate_99(G331gat,muxed95,G264gat);
xor gate_100(G332gat,muxed95,muxed37);
xor gate_101(G333gat,muxed95,G270gat);
nand gate_102(G334gat,G8gat,muxed89);
xor gate_103(G335gat,muxed95,muxed62);
nand gate_104(G336gat,muxed89,G21gat);
xor gate_105(G337gat,muxed95,G276gat);
nand gate_106(G338gat,muxed89,G34gat);
xor gate_107(G339gat,muxed95,G279gat);
nand gate_108(G340gat,muxed89,G47gat);
xor gate_109(G341gat,muxed95,G282gat);
nand gate_110(G342gat,muxed89,G60gat);
xor gate_111(G343gat,muxed95,G285gat);
nand gate_112(G344gat,muxed89,muxed26);
nand gate_113(G345gat,muxed89,G86gat);
nand gate_114(G346gat,muxed89,G99gat);
nand gate_115(G347gat,muxed89,G112gat);
nand gate_116(G348gat,muxed63,G300gat);
nand gate_117(G349gat,G331gat,muxed65);
nand gate_118(G350gat,G332gat,G302gat);
nand gate_119(G351gat,G333gat,muxed10);
nand gate_120(G352gat,muxed60,G304gat);
nand gate_121(G353gat,G337gat,G305gat);
nand gate_122(G354gat,muxed42,G306gat);
nand gate_123(G355gat,G341gat,G307gat);
nand gate_124(G356gat,G343gat,G308gat);
and gate_125(G357gat,muxed74,muxed64,G350gat,muxed8,muxed58,G353gat,muxed41,muxed24,G356gat);
not gate_126(G360gat,muxed55);
not gate_127(G370gat,muxed55);
nand gate_128(G371gat,G14gat,muxed52);
nand gate_129(G372gat,muxed52,G27gat);
nand gate_130(G373gat,muxed52,G40gat);
nand gate_131(G374gat,muxed52,G53gat);
nand gate_132(G375gat,muxed52,G66gat);
nand gate_133(G376gat,muxed52,G79gat);
nand gate_134(G377gat,muxed52,G92gat);
nand gate_135(G378gat,muxed52,G105gat);
nand gate_136(G379gat,muxed52,G115gat);
nand gate_137(G380gat,G4gat,G242gat,G334gat,G371gat);
nand gate_138(G381gat,muxed61,G336gat,G372gat,muxed76);
nand gate_139(G386gat,muxed36,G338gat,G373gat,G30gat);
nand gate_140(G393gat,G254gat,G340gat,muxed59,G43gat);
nand gate_141(G399gat,muxed28,muxed98,G375gat,G56gat);
nand gate_142(G404gat,G256gat,muxed83,G376gat,G69gat);
nand gate_143(G407gat,G257gat,G345gat,G377gat,G82gat);
nand gate_144(G411gat,G258gat,G346gat,G378gat,G95gat);
nand gate_145(G414gat,G259gat,G347gat,muxed4,G108gat);
not gate_146(G415gat,G380gat);
and gate_147(G416gat,G381gat,muxed30,G393gat,muxed25,muxed82,G407gat,G411gat,muxed2);
not gate_148(G417gat,G393gat);
not gate_149(G418gat,muxed82);
not gate_150(G419gat,G407gat);
not gate_151(G420gat,G411gat);
nor gate_152(G421gat,G415gat,muxed101);
nand gate_153(G422gat,muxed30,G417gat);
nand gate_154(G425gat,muxed30,G393gat,muxed80,muxed25);
nand gate_155(G428gat,muxed25,G393gat,G419gat);
nand gate_156(G429gat,muxed30,G393gat,G407gat,G420gat);
nand gate_157(G430gat,G381gat,muxed30,G422gat,muxed25);
nand gate_158(G431gat,G381gat,muxed30,muxed77,G428gat);
nand gate_159(G432gat,G381gat,G422gat,muxed77,muxed75);
assign muxed0 = keyinput0 ? G233gat : muxed101;
assign muxed1 = keyinput1 ? muxed23 : G381gat;
assign muxed2 = keyinput2 ? G414gat : G263gat;
assign muxed3 = keyinput3 ? G159gat : G414gat;
assign muxed4 = keyinput4 ? muxed91 : G258gat;
assign muxed5 = keyinput5 ? muxed100 : muxed91;
assign muxed6 = keyinput6 ? muxed53 : muxed46;
assign muxed7 = keyinput7 ? muxed56 : G304gat;
assign muxed8 = keyinput8 ? muxed32 : G343gat;
assign muxed9 = keyinput9 ? muxed33 : muxed32;
assign muxed10 = keyinput10 ? muxed44 : G306gat;
assign muxed11 = keyinput11 ? G339gat : muxed44;
assign muxed12 = keyinput12 ? muxed20 : muxed47;
assign muxed13 = keyinput13 ? G250gat : muxed20;
assign muxed14 = keyinput14 ? G255gat : muxed30;
assign muxed15 = keyinput15 ? muxed31 : G143gat;
assign muxed16 = keyinput16 ? muxed35 : G203gat;
assign muxed17 = keyinput17 ? muxed78 : muxed35;
assign muxed18 = keyinput18 ? muxed13 : muxed38;
assign muxed19 = keyinput19 ? G188gat : muxed13;
assign muxed20 = keyinput20 ? G290gat : G150gat;
assign muxed21 = keyinput21 ? muxed0 : G356gat;
assign muxed22 = keyinput22 ? muxed1 : G168gat;
assign muxed23 = keyinput23 ? muxed54 : muxed41;
assign muxed24 = keyinput24 ? G355gat : muxed54;
assign muxed25 = keyinput25 ? muxed93 : G150gat;
assign muxed26 = keyinput26 ? G73gat : muxed93;
assign muxed27 = keyinput27 ? muxed96 : muxed41;
assign muxed28 = keyinput28 ? muxed14 : G168gat;
assign muxed29 = keyinput29 ? G195gat : muxed14;
assign muxed30 = keyinput30 ? muxed15 : G380gat;
assign muxed31 = keyinput31 ? muxed9 : muxed32;
assign muxed32 = keyinput32 ? G351gat : muxed9;
assign muxed33 = keyinput33 ? muxed16 : G260gat;
assign muxed34 = keyinput34 ? muxed69 : muxed16;
assign muxed35 = keyinput35 ? G386gat : muxed21;
assign muxed36 = keyinput36 ? muxed18 : G165gat;
assign muxed37 = keyinput37 ? muxed66 : muxed18;
assign muxed38 = keyinput38 ? G191gat : G239gat;
assign muxed39 = keyinput39 ? G142gat : muxed93;
assign muxed40 = keyinput40 ? muxed94 : G190gat;
assign muxed41 = keyinput41 ? G354gat : G260gat;
assign muxed42 = keyinput42 ? muxed11 : G197gat;
assign muxed43 = keyinput43 ? G180gat : muxed11;
assign muxed44 = keyinput44 ? G303gat : G191gat;
assign muxed45 = keyinput45 ? muxed12 : muxed31;
assign muxed46 = keyinput46 ? G171gat : muxed12;
assign muxed47 = keyinput47 ? G293gat : G353gat;
assign muxed48 = keyinput48 ? G243gat : G183gat;
assign muxed49 = keyinput49 ? G174gat : G254gat;
assign muxed50 = keyinput50 ? G236gat : muxed91;
assign muxed51 = keyinput51 ? G379gat : muxed92;
assign muxed52 = keyinput52 ? muxed6 : muxed29;
assign muxed53 = keyinput53 ? G360gat : muxed1;
assign muxed54 = keyinput54 ? G416gat : G360gat;
assign muxed55 = keyinput55 ? muxed7 : G386gat;
assign muxed56 = keyinput56 ? muxed73 : G185gat;
assign muxed57 = keyinput57 ? muxed3 : muxed73;
assign muxed58 = keyinput58 ? G352gat : G180gat;
assign muxed59 = keyinput59 ? G374gat : G352gat;
assign muxed60 = keyinput60 ? G335gat : G255gat;
assign muxed61 = keyinput61 ? muxed99 : G335gat;
assign muxed62 = keyinput62 ? G273gat : muxed35;
assign muxed63 = keyinput63 ? G330gat : muxed64;
assign muxed64 = keyinput64 ? G349gat : G428gat;
assign muxed65 = keyinput65 ? G301gat : G257gat;
assign muxed66 = keyinput66 ? G267gat : G301gat;
assign muxed67 = keyinput67 ? muxed34 : G250gat;
assign muxed68 = keyinput68 ? G294gat : muxed34;
assign muxed69 = keyinput69 ? muxed85 : G303gat;
assign muxed70 = keyinput70 ? muxed81 : muxed85;
assign muxed71 = keyinput71 ? G227gat : muxed10;
assign muxed72 = keyinput72 ? muxed57 : muxed25;
assign muxed73 = keyinput73 ? G357gat : G416gat;
assign muxed74 = keyinput74 ? G348gat : muxed48;
assign muxed75 = keyinput75 ? G429gat : G348gat;
assign muxed76 = keyinput76 ? G17gat : muxed77;
assign muxed77 = keyinput77 ? muxed17 : muxed44;
assign muxed78 = keyinput78 ? G425gat : muxed38;
assign muxed79 = keyinput79 ? G130gat : G425gat;
assign muxed80 = keyinput80 ? G418gat : G138gat;
assign muxed81 = keyinput81 ? G344gat : G418gat;
assign muxed82 = keyinput82 ? G404gat : G157gat;
assign muxed83 = keyinput83 ? muxed70 : G157gat;
assign muxed84 = keyinput84 ? G192gat : muxed70;
assign muxed85 = keyinput85 ? G288gat : G336gat;
assign muxed86 = keyinput86 ? G184gat : G171gat;
assign muxed87 = keyinput87 ? G134gat : G184gat;
assign muxed88 = keyinput88 ? G123gat : G293gat;
assign muxed89 = keyinput89 ? G319gat : muxed90;
assign muxed90 = keyinput90 ? muxed50 : G165gat;
assign muxed91 = keyinput91 ? muxed51 : G351gat;
assign muxed92 = keyinput92 ? muxed97 : muxed23;
assign muxed93 = keyinput93 ? muxed40 : G418gat;
assign muxed94 = keyinput94 ? muxed27 : muxed3;
assign muxed95 = keyinput95 ? G309gat : muxed27;
assign muxed96 = keyinput96 ? G399gat : G414gat;
assign muxed97 = keyinput97 ? muxed39 : G399gat;
assign muxed98 = keyinput98 ? muxed5 : G247gat;
assign muxed99 = keyinput99 ? G246gat : muxed5;
assign muxed100 = keyinput100 ? G342gat : G250gat;
assign muxed101 = keyinput101 ? muxed22 : G342gat;
endmodule
