`timescale 1ns / 1ps
// Verilog
// c499
// Ninputs 41
// Noutputs 32
// NtotalGates 202
// XOR2 104
// AND2 40
// NOT1 40
// AND4 8
// OR4 2
// AND5 8

module top (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
                  N753,N754,N755,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
                  keyinput60, keyinput61, keyinput62, keyinput63,
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
        keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
        keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
        keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
        keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
        keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
        keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
        keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
                  keyinput144, keyinput145,
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150,
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155,
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160,
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165,
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170,
        keyinput171, keyinput172, keyinput173, keyinput174, keyinput175,
        keyinput176, keyinput177, keyinput178, keyinput179, keyinput180,
        keyinput181, keyinput182, keyinput183, keyinput184, keyinput185,
        keyinput186);

  input keyinput146, keyinput147, keyinput148, keyinput149, keyinput150;
  input keyinput151, keyinput152, keyinput153, keyinput154, keyinput155;
  input keyinput156, keyinput157, keyinput158, keyinput159, keyinput160;
  input keyinput161, keyinput162, keyinput163, keyinput164, keyinput165;
  input keyinput166, keyinput167, keyinput168, keyinput169, keyinput170;
  input keyinput171, keyinput172, keyinput173, keyinput174, keyinput175;
  input keyinput176, keyinput177, keyinput178, keyinput179, keyinput180;
  input keyinput181, keyinput182, keyinput183, keyinput184, keyinput185;
  input keyinput186;


  input keyinput64, keyinput65, keyinput66, keyinput67, keyinput68;
  input keyinput69, keyinput70, keyinput71, keyinput72, keyinput73;
  input keyinput74, keyinput75, keyinput76, keyinput77, keyinput78;
  input keyinput79, keyinput80, keyinput81, keyinput82, keyinput83;
  input keyinput84, keyinput85, keyinput86, keyinput87, keyinput88;
  input keyinput89, keyinput90, keyinput91, keyinput92, keyinput93;
  input keyinput94, keyinput95, keyinput96, keyinput97, keyinput98;
  input keyinput99, keyinput100, keyinput101, keyinput102, keyinput103;
  input keyinput104, keyinput105, keyinput106, keyinput107, keyinput108;
  input keyinput109, keyinput110, keyinput111, keyinput112, keyinput113;
  input keyinput114, keyinput115, keyinput116, keyinput117, keyinput118;
  input keyinput119, keyinput120, keyinput121, keyinput122, keyinput123;
  input keyinput124, keyinput125, keyinput126, keyinput127, keyinput128;
  input keyinput129, keyinput130, keyinput131, keyinput132, keyinput133;
  input keyinput134, keyinput135, keyinput136, keyinput137, keyinput138;
  input keyinput139, keyinput140, keyinput141, keyinput142, keyinput143;
  input keyinput144, keyinput145;

  wire KeyWire_0_1 , KeyWire_0_2;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31, keyinput32, keyinput33, keyinput34;
  input keyinput35, keyinput36, keyinput37, keyinput38, keyinput39;
  input keyinput40, keyinput41, keyinput42, keyinput43, keyinput44;
  input keyinput45, keyinput46, keyinput47, keyinput48, keyinput49;
  input keyinput50, keyinput51, keyinput52, keyinput53, keyinput54;
  input keyinput55, keyinput56, keyinput57, keyinput58, keyinput59;
  input keyinput60, keyinput61, keyinput62, keyinput63;

  wire [0:63] keyinput_Wire_0;
  wire [0:32] KeyNOTWire_0;

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;

output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723;

  xor XOR2_1 (keyinput_Wire_0[0], N1, N5);
  xor keyGate_0_0(KeyNOTWire_0[0], keyinput0, keyinput_Wire_0[0]);
  not KeyNOTGate_0_0(N250, KeyNOTWire_0[0]);
  xor XOR2_2 (keyinput_Wire_0[1], N9, N13);
  xnor keyGate_0_1(KeyNOTWire_0[1], keyinput1, keyinput_Wire_0[1]);
  not KeyNOTGate_0_1(N251, KeyNOTWire_0[1]);
  xor XOR2_3 (keyinput_Wire_0[2], N17, N21);
  xor keyGate_0_2(N252, keyinput2, keyinput_Wire_0[2]);
  xor XOR2_4 (keyinput_Wire_0[3], N25, N29);
  xor keyGate_0_3(KeyNOTWire_0[2], keyinput3, keyinput_Wire_0[3]);
  not KeyNOTGate_0_2(N253, KeyNOTWire_0[2]);
  xor XOR2_5 (keyinput_Wire_0[4], N33, N37);
  xor keyGate_0_4(KeyNOTWire_0[3], keyinput4, keyinput_Wire_0[4]);
  not KeyNOTGate_0_3(N254, KeyNOTWire_0[3]);
  xor XOR2_6 (keyinput_Wire_0[5], N41, N45);
  xnor keyGate_0_5(N255, keyinput5, keyinput_Wire_0[5]);
  xor XOR2_7 (keyinput_Wire_0[6], N49, N53);
  xor keyGate_0_6(N256, keyinput6, keyinput_Wire_0[6]);
  xor XOR2_8 (keyinput_Wire_0[7], N57, N61);
  xor keyGate_0_7(N257, keyinput7, keyinput_Wire_0[7]);
  xor XOR2_9 (keyinput_Wire_0[8], N65, N69);
  xnor keyGate_0_8(KeyNOTWire_0[4], keyinput8, keyinput_Wire_0[8]);
  not KeyNOTGate_0_4(N258, KeyNOTWire_0[4]);
xor XOR2_10 (N259, N73, N77);
xor XOR2_11 (N260, N81, N85);
xor XOR2_12 (N261, N89, N93);
xor XOR2_13 (N262, N97, N101);
xor XOR2_14 (N263, N105, N109);
xor XOR2_15 (N264, N113, N117);
xor XOR2_16 (N265, N121, N125);
and AND2_17 (N266, N129, N137);
and AND2_18 (N267, N130, N137);
and AND2_19 (N268, N131, N137);
and AND2_20 (N269, N132, N137);
and AND2_21 (N270, N133, N137);
and AND2_22 (N271, N134, N137);
and AND2_23 (N272, N135, N137);
and AND2_24 (N273, N136, N137);
xor XOR2_25 (N274, N1, N17);
xor XOR2_26 (N275, N33, N49);
xor XOR2_27 (N276, N5, N21);
xor XOR2_28 (N277, N37, N53);
xor XOR2_29 (N278, N9, N25);
xor XOR2_30 (N279, N41, N57);
xor XOR2_31 (N280, N13, N29);
xor XOR2_32 (N281, N45, N61);
xor XOR2_33 (N282, N65, N81);
xor XOR2_34 (N283, N97, N113);
xor XOR2_35 (N284, N69, N85);
xor XOR2_36 (N285, N101, N117);
xor XOR2_37 (N286, N73, N89);
xor XOR2_38 (N287, N105, N121);
xor XOR2_39 (N288, N77, N93);
xor XOR2_40 (N289, N109, N125);
  xor XOR2_41 (keyinput_Wire_0[9], N250, N251);
  xor keyGate_0_9(KeyNOTWire_0[5], keyinput9, keyinput_Wire_0[9]);
  not KeyNOTGate_0_5(N290, KeyNOTWire_0[5]);
  xor XOR2_42 (keyinput_Wire_0[10], N252, N253);
  xnor keyGate_0_10(KeyNOTWire_0[6], keyinput10, keyinput_Wire_0[10]);
  not KeyNOTGate_0_6(N293, KeyNOTWire_0[6]);
  xor XOR2_43 (keyinput_Wire_0[11], N254, N255);
  xnor keyGate_0_11(N296, keyinput11, keyinput_Wire_0[11]);
  xor XOR2_44 (keyinput_Wire_0[12], N256, N257);
  xnor keyGate_0_12(KeyNOTWire_0[7], keyinput12, keyinput_Wire_0[12]);
  not KeyNOTGate_0_7(N299, KeyNOTWire_0[7]);
  xor XOR2_45 (keyinput_Wire_0[13], N258, N259);
  xor keyGate_0_13(KeyNOTWire_0[8], keyinput13, keyinput_Wire_0[13]);
  not KeyNOTGate_0_8(N302, KeyNOTWire_0[8]);
  xor XOR2_46 (keyinput_Wire_0[14], N260, N261);
  xor keyGate_0_14(KeyNOTWire_0[9], keyinput14, keyinput_Wire_0[14]);
  not KeyNOTGate_0_9(N305, KeyNOTWire_0[9]);
  xor XOR2_47 (keyinput_Wire_0[15], N262, N263);
  xnor keyGate_0_15(KeyNOTWire_0[10], keyinput15, keyinput_Wire_0[15]);
  not KeyNOTGate_0_10(N308, KeyNOTWire_0[10]);
  xor XOR2_48 (keyinput_Wire_0[16], N264, N265);
  xnor keyGate_0_16(KeyNOTWire_0[11], keyinput16, keyinput_Wire_0[16]);
  not KeyNOTGate_0_11(N311, KeyNOTWire_0[11]);
xor XOR2_49 (N314, N274, N275);
xor XOR2_50 (N315, N276, N277);
xor XOR2_51 (N316, N278, N279);
xor XOR2_52 (N317, N280, N281);
xor XOR2_53 (N318, N282, N283);
xor XOR2_54 (N319, N284, N285);
xor XOR2_55 (N320, N286, N287);
xor XOR2_56 (N321, N288, N289);
xor XOR2_57 (N338, N290, N293);
xor XOR2_58 (N339, N296, N299);
xor XOR2_59 (N340, N290, N296);
xor XOR2_60 (N341, N293, N299);
xor XOR2_61 (N342, N302, N305);
xor XOR2_62 (N343, N308, N311);
xor XOR2_63 (N344, N302, N308);
xor XOR2_64 (N345, N305, N311);
xor XOR2_65 (N346, N266, N342);
xor XOR2_66 (N347, N267, N343);
xor XOR2_67 (N348, N268, N344);
xor XOR2_68 (N349, N269, N345);
xor XOR2_69 (N350, N270, N338);
xor XOR2_70 (N351, N271, N339);
xor XOR2_71 (N352, N272, N340);
xor XOR2_72 (N353, N273, N341);
xor XOR2_73 (N354, N314, N346);
xor XOR2_74 (N367, N315, N347);
xor XOR2_75 (N380, N316, N348);
xor XOR2_76 (N393, N317, N349);
xor XOR2_77 (N406, N318, N350);
xor XOR2_78 (N419, N319, N351);
xor XOR2_79 (N432, N320, N352);
xor XOR2_80 (N445, N321, N353);
not NOT1_81 (N554, N354);
not NOT1_82 (N555, N367);
not NOT1_83 (N556, N380);
not NOT1_84 (N557, N354);
not NOT1_85 (N558, N367);
not NOT1_86 (N559, N393);
not NOT1_87 (N560, N354);
not NOT1_88 (N561, N380);
not NOT1_89 (N562, N393);
not NOT1_90 (N563, N367);
not NOT1_91 (N564, N380);
not NOT1_92 (N565, N393);
not NOT1_93 (N566, N419);
not NOT1_94 (N567, N445);
not NOT1_95 (N568, N419);
not NOT1_96 (N569, N432);
not NOT1_97 (N570, N406);
not NOT1_98 (N571, N445);
not NOT1_99 (N572, N406);
not NOT1_100 (N573, N432);
not NOT1_101 (N574, N406);
not NOT1_102 (N575, N419);
not NOT1_103 (N576, N432);
not NOT1_104 (N577, N406);
not NOT1_105 (N578, N419);
not NOT1_106 (N579, N445);
not NOT1_107 (N580, N406);
not NOT1_108 (N581, N432);
not NOT1_109 (N582, N445);
not NOT1_110 (N583, N419);
not NOT1_111 (N584, N432);
not NOT1_112 (N585, N445);
not NOT1_113 (N586, N367);
not NOT1_114 (N587, N393);
not NOT1_115 (N588, N367);
not NOT1_116 (N589, N380);
not NOT1_117 (N590, N354);
not NOT1_118 (N591, N393);
not NOT1_119 (N592, N354);
not NOT1_120 (N593, N380);
and AND4_121 (N594, N554, N555, N556, N393);
and AND4_122 (N595, N557, N558, N380, N559);
and AND4_123 (N596, N560, N367, N561, N562);
and AND4_124 (N597, N354, N563, N564, N565);
and AND4_125 (N598, N574, N575, N576, N445);
and AND4_126 (N599, N577, N578, N432, N579);
and AND4_127 (N600, N580, N419, N581, N582);
and AND4_128 (N601, N406, N583, N584, N585);
or OR4_129 (N602, N594, N595, N596, N597);
or OR4_130 (N607, N598, N599, N600, N601);
  and AND5_131 (keyinput_Wire_0[17], N406, N566, N432, N567, N602);
  xnor keyGate_0_17(KeyNOTWire_0[12], keyinput17, keyinput_Wire_0[17]);
  not KeyNOTGate_0_12(N620, KeyNOTWire_0[12]);
  and AND5_132 (keyinput_Wire_0[18], N406, N568, N569, N445, N602);
  xnor keyGate_0_18(N625, keyinput18, keyinput_Wire_0[18]);
  and AND5_133 (keyinput_Wire_0[19], N570, N419, N432, N571, N602);
  xnor keyGate_0_19(N630, keyinput19, keyinput_Wire_0[19]);
  and AND5_134 (keyinput_Wire_0[20], N572, N419, N573, N445, N602);
  xnor keyGate_0_20(KeyNOTWire_0[13], keyinput20, keyinput_Wire_0[20]);
  not KeyNOTGate_0_13(N635, KeyNOTWire_0[13]);
  and AND5_135 (keyinput_Wire_0[21], N354, N586, N380, N587, N607);
  xor keyGate_0_21(KeyNOTWire_0[14], keyinput21, keyinput_Wire_0[21]);
  not KeyNOTGate_0_14(N640, KeyNOTWire_0[14]);
  and AND5_136 (keyinput_Wire_0[22], N354, N588, N589, N393, N607);
  xnor keyGate_0_22(KeyNOTWire_0[15], keyinput22, keyinput_Wire_0[22]);
  not KeyNOTGate_0_15(N645, KeyNOTWire_0[15]);
  and AND5_137 (keyinput_Wire_0[23], N590, N367, N380, N591, N607);
  xnor keyGate_0_23(KeyNOTWire_0[16], keyinput23, keyinput_Wire_0[23]);
  not KeyNOTGate_0_16(N650, KeyNOTWire_0[16]);
  and AND5_138 (keyinput_Wire_0[24], N592, N367, N593, N393, N607);
  xor keyGate_0_24(KeyNOTWire_0[17], keyinput24, keyinput_Wire_0[24]);
  not KeyNOTGate_0_17(N655, KeyNOTWire_0[17]);
and AND2_139 (N692, N354, N620);
and AND2_140 (N693, N367, N620);
and AND2_141 (N694, N380, N620);
and AND2_142 (N695, N393, N620);
and AND2_143 (N696, N354, N625);
  and AND2_144 (keyinput_Wire_0[25], N367, N625);
  xor keyGate_0_25(KeyNOTWire_0[18], keyinput25, keyinput_Wire_0[25]);
  not KeyNOTGate_0_18(N697, KeyNOTWire_0[18]);
  and AND2_145 (keyinput_Wire_0[26], N380, N625);
  xnor keyGate_0_26(N698, keyinput26, keyinput_Wire_0[26]);
  and AND2_146 (keyinput_Wire_0[27], N393, N625);
  xnor keyGate_0_27(KeyNOTWire_0[19], keyinput27, keyinput_Wire_0[27]);
  not KeyNOTGate_0_19(N699, KeyNOTWire_0[19]);
  and AND2_147 (keyinput_Wire_0[28], N354, N630);
  xnor keyGate_0_28(N700, keyinput28, keyinput_Wire_0[28]);
  and AND2_148 (keyinput_Wire_0[29], N367, N630);
  xnor keyGate_0_29(N701, keyinput29, keyinput_Wire_0[29]);
  and AND2_149 (keyinput_Wire_0[30], N380, N630);
  xor keyGate_0_30(N702, keyinput30, keyinput_Wire_0[30]);
  and AND2_150 (keyinput_Wire_0[31], N393, N630);
  xnor keyGate_0_31(KeyNOTWire_0[20], keyinput31, keyinput_Wire_0[31]);
  not KeyNOTGate_0_20(N703, KeyNOTWire_0[20]);
  and AND2_151 (keyinput_Wire_0[32], N354, N635);
  xnor keyGate_0_32(KeyNOTWire_0[21], keyinput32, keyinput_Wire_0[32]);
  not KeyNOTGate_0_21(N704, KeyNOTWire_0[21]);
  and AND2_152 (keyinput_Wire_0[33], N367, N635);
  xor keyGate_0_33(N705, keyinput33, keyinput_Wire_0[33]);
  and AND2_153 (keyinput_Wire_0[34], N380, N635);
  xnor keyGate_0_34(N706, keyinput34, keyinput_Wire_0[34]);
  and AND2_154 (keyinput_Wire_0[35], N393, N635);
  xor keyGate_0_35(N707, keyinput35, keyinput_Wire_0[35]);
  and AND2_155 (keyinput_Wire_0[36], N406, N640);
  xor keyGate_0_36(N708, keyinput36, keyinput_Wire_0[36]);
  and AND2_156 (keyinput_Wire_0[37], N419, N640);
  xor keyGate_0_37(N709, keyinput37, keyinput_Wire_0[37]);
  and AND2_157 (keyinput_Wire_0[38], N432, N640);
  xnor keyGate_0_38(N710, keyinput38, keyinput_Wire_0[38]);
  and AND2_158 (keyinput_Wire_0[39], N445, N640);
  xnor keyGate_0_39(N711, keyinput39, keyinput_Wire_0[39]);
  and AND2_159 (keyinput_Wire_0[40], N406, N645);
  xor keyGate_0_40(N712, keyinput40, keyinput_Wire_0[40]);
and AND2_160 (N713, N419, N645);
and AND2_161 (N714, N432, N645);
and AND2_162 (N715, N445, N645);
and AND2_163 (N716, N406, N650);
and AND2_164 (N717, N419, N650);
and AND2_165 (N718, N432, N650);
and AND2_166 (N719, N445, N650);
and AND2_167 (N720, N406, N655);
and AND2_168 (N721, N419, N655);
and AND2_169 (N722, N432, N655);
and AND2_170 (N723, N445, N655);
xor XOR2_171 (N724, N1, N692);
xor XOR2_172 (N725, N5, N693);
xor XOR2_173 (N726, N9, N694);
xor XOR2_174 (N727, N13, N695);
xor XOR2_175 (N728, N17, N696);
xor XOR2_176 (N729, N21, N697);
xor XOR2_177 (N730, N25, N698);
xor XOR2_178 (N731, N29, N699);
xor XOR2_179 (N732, N33, N700);
  xor XOR2_180 (keyinput_Wire_0[41], N37, N701);
  xnor keyGate_0_41(N733, keyinput41, keyinput_Wire_0[41]);
  xor XOR2_181 (keyinput_Wire_0[42], N41, N702);
  xor keyGate_0_42(KeyNOTWire_0[22], keyinput42, keyinput_Wire_0[42]);
  not KeyNOTGate_0_22(N734, KeyNOTWire_0[22]);
  xor XOR2_182 (keyinput_Wire_0[43], N45, N703);
  xnor keyGate_0_43(KeyNOTWire_0[23], keyinput43, keyinput_Wire_0[43]);
  not KeyNOTGate_0_23(N735, KeyNOTWire_0[23]);
  xor XOR2_183 (keyinput_Wire_0[44], N49, N704);
  xor keyGate_0_44(KeyNOTWire_0[24], keyinput44, keyinput_Wire_0[44]);
  not KeyNOTGate_0_24(N736, KeyNOTWire_0[24]);
  xor XOR2_184 (keyinput_Wire_0[45], N53, N705);
  xor keyGate_0_45(KeyNOTWire_0[25], keyinput45, keyinput_Wire_0[45]);
  not KeyNOTGate_0_25(N737, KeyNOTWire_0[25]);
  xor XOR2_185 (keyinput_Wire_0[46], N57, N706);
  xor keyGate_0_46(N738, keyinput46, keyinput_Wire_0[46]);
  xor XOR2_186 (keyinput_Wire_0[47], N61, N707);
  xnor keyGate_0_47(N739, keyinput47, keyinput_Wire_0[47]);
  xor XOR2_187 (keyinput_Wire_0[48], N65, N708);
  xnor keyGate_0_48(N740, keyinput48, keyinput_Wire_0[48]);
  xor XOR2_188 (keyinput_Wire_0[49], N69, N709);
  xor keyGate_0_49(N741, keyinput49, keyinput_Wire_0[49]);
  xor XOR2_189 (keyinput_Wire_0[50], N73, N710);
  xnor keyGate_0_50(KeyNOTWire_0[26], keyinput50, keyinput_Wire_0[50]);
  not KeyNOTGate_0_26(N742, KeyNOTWire_0[26]);
  xor XOR2_190 (keyinput_Wire_0[51], N77, N711);
  xor keyGate_0_51(KeyNOTWire_0[27], keyinput51, keyinput_Wire_0[51]);
  not KeyNOTGate_0_27(N743, KeyNOTWire_0[27]);
  xor XOR2_191 (keyinput_Wire_0[52], N81, N712);
  xor keyGate_0_52(KeyNOTWire_0[28], keyinput52, keyinput_Wire_0[52]);
  not KeyNOTGate_0_28(N744, KeyNOTWire_0[28]);
  xor XOR2_192 (keyinput_Wire_0[53], N85, N713);
  xor keyGate_0_53(N745, keyinput53, keyinput_Wire_0[53]);
  xor XOR2_193 (keyinput_Wire_0[54], N89, N714);
  xnor keyGate_0_54(KeyNOTWire_0[29], keyinput54, keyinput_Wire_0[54]);
  not KeyNOTGate_0_29(N746, KeyNOTWire_0[29]);
  xor XOR2_194 (keyinput_Wire_0[55], N93, N715);
  xor keyGate_0_55(KeyNOTWire_0[30], keyinput55, keyinput_Wire_0[55]);
  not KeyNOTGate_0_30(N747, KeyNOTWire_0[30]);
  xor XOR2_195 (keyinput_Wire_0[56], N97, N716);
  xor keyGate_0_56(N748, keyinput56, keyinput_Wire_0[56]);
  xor XOR2_196 (keyinput_Wire_0[57], N101, N717);
  xnor keyGate_0_57(KeyNOTWire_0[31], keyinput57, keyinput_Wire_0[57]);
  not KeyNOTGate_0_31(N749, KeyNOTWire_0[31]);
  xor XOR2_197 (keyinput_Wire_0[58], N105, N718);
  xor keyGate_0_58(KeyNOTWire_0[32], keyinput58, keyinput_Wire_0[58]);
  not KeyNOTGate_0_32(KeyWire_0_1, KeyNOTWire_0[32]);
  xor flip_it (N750, KeyWire_0_1, KeyWire_0_2 );
  xor XOR2_198 (keyinput_Wire_0[59], N109, N719);
  xor keyGate_0_59(N751, keyinput59, keyinput_Wire_0[59]);
  xor XOR2_199 (keyinput_Wire_0[60], N113, N720);
  xor keyGate_0_60(N752, keyinput60, keyinput_Wire_0[60]);
  xor XOR2_200 (keyinput_Wire_0[61], N117, N721);
  xnor keyGate_0_61(N753, keyinput61, keyinput_Wire_0[61]);
  xor XOR2_201 (keyinput_Wire_0[62], N121, N722);
  xor keyGate_0_62(N754, keyinput62, keyinput_Wire_0[62]);
  xor XOR2_202 (keyinput_Wire_0[63], N125, N723);
  xnor keyGate_0_63(N755, keyinput63, keyinput_Wire_0[63]);

AntiSAT some_name( KeyWire_0_2, N105, N97, N73, N101, N29, N81, N130, N17, N45, N13, N117, N9, N121, N113, N25, N33, N1, N65, N135, N61, N93, N133, N134, N89, N21, N132, N49, N109, N136, N131, N57, N137, N53, N125, N77, N85, N129, N41, N5, N37, N69, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145,
       keyinput146, keyinput147, keyinput148, keyinput149, keyinput150,
       keyinput151, keyinput152, keyinput153, keyinput154, keyinput155,
       keyinput156, keyinput157, keyinput158, keyinput159, keyinput160,
       keyinput161, keyinput162, keyinput163, keyinput164, keyinput165,
       keyinput166, keyinput167, keyinput168, keyinput169, keyinput170,
       keyinput171, keyinput172, keyinput173, keyinput174, keyinput175,
       keyinput176, keyinput177, keyinput178, keyinput179, keyinput180,
       keyinput181, keyinput182, keyinput183, keyinput184, keyinput185,
       keyinput186);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N105, N97, N73, N101, N29, N81, N130, N17, N45, N13, N117, N9, N121, N113, N25, N33, N1, N65, N135, N61, N93, N133, N134, N89, N21, N132, N49, N109, N136, N131, N57, N137, N53, N125, N77, N85, N129, N41, N5, N37, N69, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145 ,
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150,
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155,
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160,
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165,
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170,
        keyinput171, keyinput172, keyinput173, keyinput174, keyinput175,
        keyinput176, keyinput177, keyinput178, keyinput179, keyinput180,
        keyinput181, keyinput182, keyinput183, keyinput184, keyinput185,
        keyinput186);

  input keyinput146, keyinput147, keyinput148, keyinput149, keyinput150;
  input keyinput151, keyinput152, keyinput153, keyinput154, keyinput155;
  input keyinput156, keyinput157, keyinput158, keyinput159, keyinput160;
  input keyinput161, keyinput162, keyinput163, keyinput164, keyinput165;
  input keyinput166, keyinput167, keyinput168, keyinput169, keyinput170;
  input keyinput171, keyinput172, keyinput173, keyinput174, keyinput175;
  input keyinput176, keyinput177, keyinput178, keyinput179, keyinput180;
  input keyinput181, keyinput182, keyinput183, keyinput184, keyinput185;
  input keyinput186;

  wire [0:40] keyNTin_Wire_1;
  wire [0:19] KeyNOTWire_1;

  input N105, N97, N73, N101, N29, N81, N130, N17, N45, N13, N117, N9, N121, N113, N25, N33, N1, N65, N135, N61, N93, N133, N134, N89, N21, N132, N49, N109, N136, N131, N57, N137, N53, N125, N77, N85, N129, N41, N5, N37, N69;
  input keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83 ;

  xor  KeyGate0 (newWire_0, N105, keyinput64);
  xnor KeyGate1 (keyNTin_Wire_1[0], N97, keyinput65);
  xor keyNTinGate_1_0(newWire_1, keyinput146, keyNTin_Wire_1[0]);
  xor  KeyGate2 (newWire_2, N73, keyinput66);
  xor  KeyGate3 (newWire_3, N101, keyinput67);
  xor  KeyGate4 (keyNTin_Wire_1[1], N29, keyinput68);
  xor keyNTinGate_1_1(newWire_4, keyinput147, keyNTin_Wire_1[1]);
  xor  KeyGate5 (newWire_5, N81, keyinput69);
  xor  KeyGate6 (newWire_6, N130, keyinput70);
  xnor KeyGate7 (newWire_7, N17, keyinput71);
  xnor KeyGate8 (newWire_8, N45, keyinput72);
  xnor KeyGate9 (keyNTin_Wire_1[2], N13, keyinput73);
  xnor keyNTinGate_1_2(KeyNOTWire_1[0], keyinput148, keyNTin_Wire_1[2]);
  not KeyNOTGate_1_0(newWire_9, KeyNOTWire_1[0]);
  xnor KeyGate10 (keyNTin_Wire_1[3], N117, keyinput74);
  xnor keyNTinGate_1_3(KeyNOTWire_1[1], keyinput149, keyNTin_Wire_1[3]);
  not KeyNOTGate_1_1(newWire_10, KeyNOTWire_1[1]);
  xor  KeyGate11 (keyNTin_Wire_1[4], N9, keyinput75);
  xnor keyNTinGate_1_4(KeyNOTWire_1[2], keyinput150, keyNTin_Wire_1[4]);
  not KeyNOTGate_1_2(newWire_11, KeyNOTWire_1[2]);
  xor  KeyGate12 (newWire_12, N121, keyinput76);
  xor  KeyGate13 (newWire_13, N113, keyinput77);
  xor  KeyGate14 (newWire_14, N25, keyinput78);
  xor  KeyGate15 (newWire_15, N33, keyinput79);
  xnor KeyGate16 (newWire_16, N1, keyinput80);
  xnor KeyGate17 (newWire_17, N65, keyinput81);
  xnor KeyGate18 (keyNTin_Wire_1[5], N135, keyinput82);
  xnor keyNTinGate_1_5(newWire_18, keyinput151, keyNTin_Wire_1[5]);
  xor  KeyGate19 (keyNTin_Wire_1[6], N61, keyinput83);
  xor keyNTinGate_1_6(newWire_19, keyinput152, keyNTin_Wire_1[6]);
  xor  KeyGate20 (keyNTin_Wire_1[7], N93, keyinput84);
  xor keyNTinGate_1_7(newWire_20, keyinput153, keyNTin_Wire_1[7]);
  xnor KeyGate21 (newWire_21, N133, keyinput85);
  xnor KeyGate22 (newWire_22, N134, keyinput86);
  xor  KeyGate23 (keyNTin_Wire_1[8], N89, keyinput87);
  xor keyNTinGate_1_8(newWire_23, keyinput154, keyNTin_Wire_1[8]);
  xor  KeyGate24 (newWire_24, N21, keyinput88);
  xor  KeyGate25 (keyNTin_Wire_1[9], N132, keyinput89);
  xor keyNTinGate_1_9(newWire_25, keyinput155, keyNTin_Wire_1[9]);
  xor  KeyGate26 (keyNTin_Wire_1[10], N49, keyinput90);
  xnor keyNTinGate_1_10(KeyNOTWire_1[3], keyinput156, keyNTin_Wire_1[10]);
  not KeyNOTGate_1_3(newWire_26, KeyNOTWire_1[3]);
  xor  KeyGate27 (keyNTin_Wire_1[11], N109, keyinput91);
  xor keyNTinGate_1_11(KeyNOTWire_1[4], keyinput157, keyNTin_Wire_1[11]);
  not KeyNOTGate_1_4(newWire_27, KeyNOTWire_1[4]);
  xor  KeyGate28 (newWire_28, N136, keyinput92);
  xnor KeyGate29 (keyNTin_Wire_1[12], N131, keyinput93);
  xnor keyNTinGate_1_12(newWire_29, keyinput158, keyNTin_Wire_1[12]);
  xor  KeyGate30 (newWire_30, N57, keyinput94);
  xnor KeyGate31 (keyNTin_Wire_1[13], N137, keyinput95);
  xor keyNTinGate_1_13(newWire_31, keyinput159, keyNTin_Wire_1[13]);
  xnor KeyGate32 (newWire_32, N53, keyinput96);
  xor  KeyGate33 (newWire_33, N125, keyinput97);
  xnor KeyGate34 (newWire_34, N77, keyinput98);
  xnor KeyGate35 (newWire_35, N85, keyinput99);
  xnor KeyGate36 (keyNTin_Wire_1[14], N129, keyinput100);
  xnor keyNTinGate_1_14(KeyNOTWire_1[5], keyinput160, keyNTin_Wire_1[14]);
  not KeyNOTGate_1_5(newWire_36, KeyNOTWire_1[5]);
  xor  KeyGate37 (keyNTin_Wire_1[15], N41, keyinput101);
  xnor keyNTinGate_1_15(newWire_37, keyinput161, keyNTin_Wire_1[15]);
  xor  KeyGate38 (keyNTin_Wire_1[16], N5, keyinput102);
  xor keyNTinGate_1_16(KeyNOTWire_1[6], keyinput162, keyNTin_Wire_1[16]);
  not KeyNOTGate_1_6(newWire_38, KeyNOTWire_1[6]);
  xor  KeyGate39 (keyNTin_Wire_1[17], N37, keyinput103);
  xnor keyNTinGate_1_17(KeyNOTWire_1[7], keyinput163, keyNTin_Wire_1[17]);
  not KeyNOTGate_1_7(newWire_39, KeyNOTWire_1[7]);
  xnor KeyGate40 (newWire_40, N69, keyinput104);
  xor  KeyGate41 (newWire_41, N105, keyinput105);
  xnor KeyGate42 (newWire_42, N97, keyinput106);
  xnor KeyGate43 (keyNTin_Wire_1[18], N73, keyinput107);
  xnor keyNTinGate_1_18(KeyNOTWire_1[8], keyinput164, keyNTin_Wire_1[18]);
  not KeyNOTGate_1_8(newWire_43, KeyNOTWire_1[8]);
  xnor KeyGate44 (newWire_44, N101, keyinput108);
  xor  KeyGate45 (keyNTin_Wire_1[19], N29, keyinput109);
  xor keyNTinGate_1_19(newWire_45, keyinput165, keyNTin_Wire_1[19]);
  xnor KeyGate46 (keyNTin_Wire_1[20], N81, keyinput110);
  xor keyNTinGate_1_20(KeyNOTWire_1[9], keyinput166, keyNTin_Wire_1[20]);
  not KeyNOTGate_1_9(newWire_46, KeyNOTWire_1[9]);
  xor  KeyGate47 (keyNTin_Wire_1[21], N130, keyinput111);
  xor keyNTinGate_1_21(newWire_47, keyinput167, keyNTin_Wire_1[21]);
  xor  KeyGate48 (keyNTin_Wire_1[22], N17, keyinput112);
  xor keyNTinGate_1_22(KeyNOTWire_1[10], keyinput168, keyNTin_Wire_1[22]);
  not KeyNOTGate_1_10(newWire_48, KeyNOTWire_1[10]);
  xor  KeyGate49 (newWire_49, N45, keyinput113);
  xnor KeyGate50 (keyNTin_Wire_1[23], N13, keyinput114);
  xor keyNTinGate_1_23(newWire_50, keyinput169, keyNTin_Wire_1[23]);
  xor  KeyGate51 (newWire_51, N117, keyinput115);
  xor  KeyGate52 (newWire_52, N9, keyinput116);
  xor  KeyGate53 (newWire_53, N121, keyinput117);
  xnor KeyGate54 (newWire_54, N113, keyinput118);
  xor  KeyGate55 (keyNTin_Wire_1[24], N25, keyinput119);
  xor keyNTinGate_1_24(KeyNOTWire_1[11], keyinput170, keyNTin_Wire_1[24]);
  not KeyNOTGate_1_11(newWire_55, KeyNOTWire_1[11]);
  xor  KeyGate56 (keyNTin_Wire_1[25], N33, keyinput120);
  xor keyNTinGate_1_25(KeyNOTWire_1[12], keyinput171, keyNTin_Wire_1[25]);
  not KeyNOTGate_1_12(newWire_56, KeyNOTWire_1[12]);
  xor  KeyGate57 (newWire_57, N1, keyinput121);
  xor  KeyGate58 (keyNTin_Wire_1[26], N65, keyinput122);
  xnor keyNTinGate_1_26(KeyNOTWire_1[13], keyinput172, keyNTin_Wire_1[26]);
  not KeyNOTGate_1_13(newWire_58, KeyNOTWire_1[13]);
  xnor KeyGate59 (keyNTin_Wire_1[27], N135, keyinput123);
  xnor keyNTinGate_1_27(newWire_59, keyinput173, keyNTin_Wire_1[27]);
  xor  KeyGate60 (newWire_60, N61, keyinput124);
  xnor KeyGate61 (newWire_61, N93, keyinput125);
  xnor KeyGate62 (newWire_62, N133, keyinput126);
  xnor KeyGate63 (keyNTin_Wire_1[28], N134, keyinput127);
  xor keyNTinGate_1_28(newWire_63, keyinput174, keyNTin_Wire_1[28]);
  xnor KeyGate64 (keyNTin_Wire_1[29], N89, keyinput128);
  xor keyNTinGate_1_29(KeyNOTWire_1[14], keyinput175, keyNTin_Wire_1[29]);
  not KeyNOTGate_1_14(newWire_64, KeyNOTWire_1[14]);
  xor  KeyGate65 (keyNTin_Wire_1[30], N21, keyinput129);
  xor keyNTinGate_1_30(newWire_65, keyinput176, keyNTin_Wire_1[30]);
  xor  KeyGate66 (keyNTin_Wire_1[31], N132, keyinput130);
  xor keyNTinGate_1_31(KeyNOTWire_1[15], keyinput177, keyNTin_Wire_1[31]);
  not KeyNOTGate_1_15(newWire_66, KeyNOTWire_1[15]);
  xor  KeyGate67 (newWire_67, N49, keyinput131);
  xor  KeyGate68 (keyNTin_Wire_1[32], N109, keyinput132);
  xor keyNTinGate_1_32(newWire_68, keyinput178, keyNTin_Wire_1[32]);
  xor  KeyGate69 (keyNTin_Wire_1[33], N136, keyinput133);
  xor keyNTinGate_1_33(KeyNOTWire_1[16], keyinput179, keyNTin_Wire_1[33]);
  not KeyNOTGate_1_16(newWire_69, KeyNOTWire_1[16]);
  xnor KeyGate70 (keyNTin_Wire_1[34], N131, keyinput134);
  xor keyNTinGate_1_34(KeyNOTWire_1[17], keyinput180, keyNTin_Wire_1[34]);
  not KeyNOTGate_1_17(newWire_70, KeyNOTWire_1[17]);
  xnor KeyGate71 (newWire_71, N57, keyinput135);
  xor  KeyGate72 (newWire_72, N137, keyinput136);
  xor  KeyGate73 (newWire_73, N53, keyinput137);
  xnor KeyGate74 (keyNTin_Wire_1[35], N125, keyinput138);
  xnor keyNTinGate_1_35(newWire_74, keyinput181, keyNTin_Wire_1[35]);
  xor  KeyGate75 (newWire_75, N77, keyinput139);
  xnor KeyGate76 (keyNTin_Wire_1[36], N85, keyinput140);
  xnor keyNTinGate_1_36(newWire_76, keyinput182, keyNTin_Wire_1[36]);
  xor  KeyGate77 (newWire_77, N129, keyinput141);
  xor  KeyGate78 (keyNTin_Wire_1[37], N41, keyinput142);
  xnor keyNTinGate_1_37(newWire_78, keyinput183, keyNTin_Wire_1[37]);
  xor  KeyGate79 (keyNTin_Wire_1[38], N5, keyinput143);
  xor keyNTinGate_1_38(KeyNOTWire_1[18], keyinput184, keyNTin_Wire_1[38]);
  not KeyNOTGate_1_18(newWire_79, KeyNOTWire_1[18]);
  xor  KeyGate80 (keyNTin_Wire_1[39], N37, keyinput144);
  xor keyNTinGate_1_39(KeyNOTWire_1[19], keyinput185, keyNTin_Wire_1[39]);
  not KeyNOTGate_1_19(newWire_80, KeyNOTWire_1[19]);
  xnor KeyGate81 (newWire_81, N69, keyinput145);
  and some_function (newWire_82, newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40 );
  nand compl_function (keyNTin_Wire_1[40], newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81);
  xor keyNTinGate_1_40(newWire_83, keyinput186, keyNTin_Wire_1[40]);
  and finalAND (KeyWire_0_2, newWire_82, newWire_83);

endmodule /* AntiSAT */
