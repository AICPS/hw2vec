`timescale 1ns / 1ps
// Verilog
// c880
// Ninputs 60
// Noutputs 26
// NtotalGates 383
// NAND4 13
// AND3 12
// NAND2 60
// NAND3 14
// AND2 105
// OR2 29
// NOT1 63
// NOR2 61
// BUFF1 26

module top (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
                  N865,N866,N874,N878,N879,N880,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
                  keyinput60, keyinput61, keyinput62, keyinput63,
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
        keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
        keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
        keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
        keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
        keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
        keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
        keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
        keyinput144, keyinput145, keyinput146, keyinput147, keyinput148,
        keyinput149, keyinput150, keyinput151, keyinput152, keyinput153,
        keyinput154, keyinput155, keyinput156, keyinput157, keyinput158,
        keyinput159, keyinput160, keyinput161, keyinput162, keyinput163,
        keyinput164, keyinput165, keyinput166, keyinput167, keyinput168,
        keyinput169, keyinput170, keyinput171, keyinput172, keyinput173,
        keyinput174, keyinput175, keyinput176, keyinput177, keyinput178,
                  keyinput179, keyinput180, keyinput181, keyinput182, keyinput183,
        keyinput184, keyinput185, keyinput186, keyinput187, keyinput188,
        keyinput189, keyinput190, keyinput191, keyinput192, keyinput193,
        keyinput194, keyinput195, keyinput196, keyinput197, keyinput198,
        keyinput199, keyinput200, keyinput201, keyinput202, keyinput203,
        keyinput204, keyinput205, keyinput206, keyinput207, keyinput208,
        keyinput209, keyinput210, keyinput211, keyinput212, keyinput213,
        keyinput214, keyinput215, keyinput216, keyinput217, keyinput218,
        keyinput219, keyinput220, keyinput221, keyinput222, keyinput223,
        keyinput224, keyinput225, keyinput226, keyinput227, keyinput228,
        keyinput229, keyinput230, keyinput231, keyinput232, keyinput233,
        keyinput234, keyinput235, keyinput236, keyinput237, keyinput238,
        keyinput239, keyinput240, keyinput241, keyinput242, keyinput243);

  input keyinput184, keyinput185, keyinput186, keyinput187, keyinput188;
  input keyinput189, keyinput190, keyinput191, keyinput192, keyinput193;
  input keyinput194, keyinput195, keyinput196, keyinput197, keyinput198;
  input keyinput199, keyinput200, keyinput201, keyinput202, keyinput203;
  input keyinput204, keyinput205, keyinput206, keyinput207, keyinput208;
  input keyinput209, keyinput210, keyinput211, keyinput212, keyinput213;
  input keyinput214, keyinput215, keyinput216, keyinput217, keyinput218;
  input keyinput219, keyinput220, keyinput221, keyinput222, keyinput223;
  input keyinput224, keyinput225, keyinput226, keyinput227, keyinput228;
  input keyinput229, keyinput230, keyinput231, keyinput232, keyinput233;
  input keyinput234, keyinput235, keyinput236, keyinput237, keyinput238;
  input keyinput239, keyinput240, keyinput241, keyinput242, keyinput243;


  input keyinput64, keyinput65, keyinput66, keyinput67, keyinput68;
  input keyinput69, keyinput70, keyinput71, keyinput72, keyinput73;
  input keyinput74, keyinput75, keyinput76, keyinput77, keyinput78;
  input keyinput79, keyinput80, keyinput81, keyinput82, keyinput83;
  input keyinput84, keyinput85, keyinput86, keyinput87, keyinput88;
  input keyinput89, keyinput90, keyinput91, keyinput92, keyinput93;
  input keyinput94, keyinput95, keyinput96, keyinput97, keyinput98;
  input keyinput99, keyinput100, keyinput101, keyinput102, keyinput103;
  input keyinput104, keyinput105, keyinput106, keyinput107, keyinput108;
  input keyinput109, keyinput110, keyinput111, keyinput112, keyinput113;
  input keyinput114, keyinput115, keyinput116, keyinput117, keyinput118;
  input keyinput119, keyinput120, keyinput121, keyinput122, keyinput123;
  input keyinput124, keyinput125, keyinput126, keyinput127, keyinput128;
  input keyinput129, keyinput130, keyinput131, keyinput132, keyinput133;
  input keyinput134, keyinput135, keyinput136, keyinput137, keyinput138;
  input keyinput139, keyinput140, keyinput141, keyinput142, keyinput143;
  input keyinput144, keyinput145, keyinput146, keyinput147, keyinput148;
  input keyinput149, keyinput150, keyinput151, keyinput152, keyinput153;
  input keyinput154, keyinput155, keyinput156, keyinput157, keyinput158;
  input keyinput159, keyinput160, keyinput161, keyinput162, keyinput163;
  input keyinput164, keyinput165, keyinput166, keyinput167, keyinput168;
  input keyinput169, keyinput170, keyinput171, keyinput172, keyinput173;
  input keyinput174, keyinput175, keyinput176, keyinput177, keyinput178;
  input keyinput179, keyinput180, keyinput181, keyinput182, keyinput183;

  wire KeyWire_0_1 , KeyWire_0_2, keyinput_Wire_1;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31, keyinput32, keyinput33, keyinput34;
  input keyinput35, keyinput36, keyinput37, keyinput38, keyinput39;
  input keyinput40, keyinput41, keyinput42, keyinput43, keyinput44;
  input keyinput45, keyinput46, keyinput47, keyinput48, keyinput49;
  input keyinput50, keyinput51, keyinput52, keyinput53, keyinput54;
  input keyinput55, keyinput56, keyinput57, keyinput58, keyinput59;
  input keyinput60, keyinput61, keyinput62, keyinput63;

  wire [0:63] keyinput_Wire_0;
  wire [0:28] KeyNOTWire_0;

input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;

output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;

wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877;

nand NAND4_1 (N269, N1, N8, N13, N17);
nand NAND4_2 (N270, N1, N26, N13, N17);
and AND3_3 (N273, N29, N36, N42);
  and AND3_4 (keyinput_Wire_0[0], N1, N26, N51);
  xor keyGate_0_0(N276, keyinput0, keyinput_Wire_0[0]);
  nand NAND4_5 (keyinput_Wire_0[1], N1, N8, N51, N17);
  xnor keyGate_0_1(KeyNOTWire_0[0], keyinput1, keyinput_Wire_0[1]);
  not KeyNOTGate_0_0(N279, KeyNOTWire_0[0]);
nand NAND4_6 (N280, N1, N8, N13, N55);
nand NAND4_7 (N284, N59, N42, N68, N72);
nand NAND2_8 (N285, N29, N68);
nand NAND3_9 (N286, N59, N68, N74);
  and AND3_10 (keyinput_Wire_0[2], N29, N75, N80);
  xnor keyGate_0_2(KeyNOTWire_0[1], keyinput2, keyinput_Wire_0[2]);
  not KeyNOTGate_0_1(N287, KeyNOTWire_0[1]);
and AND3_11 (N290, N29, N75, N42);
and AND3_12 (N291, N29, N36, N80);
and AND3_13 (N292, N29, N36, N42);
and AND3_14 (N293, N59, N75, N80);
  and AND3_15 (keyinput_Wire_0[3], N59, N75, N42);
  xnor keyGate_0_3(N294, keyinput3, keyinput_Wire_0[3]);
and AND3_16 (N295, N59, N36, N80);
and AND3_17 (N296, N59, N36, N42);
and AND2_18 (N297, N85, N86);
or OR2_19 (N298, N87, N88);
nand NAND2_20 (N301, N91, N96);
or OR2_21 (N302, N91, N96);
nand NAND2_22 (N303, N101, N106);
or OR2_23 (N304, N101, N106);
nand NAND2_24 (N305, N111, N116);
or OR2_25 (N306, N111, N116);
nand NAND2_26 (N307, N121, N126);
or OR2_27 (N308, N121, N126);
and AND2_28 (N309, N8, N138);
  not NOT1_29 (keyinput_Wire_0[4], N268);
  xnor keyGate_0_4(KeyNOTWire_0[2], keyinput4, keyinput_Wire_0[4]);
  not KeyNOTGate_0_2(N310, KeyNOTWire_0[2]);
and AND2_30 (N316, N51, N138);
and AND2_31 (N317, N17, N138);
and AND2_32 (N318, N152, N138);
  nand NAND2_33 (keyinput_Wire_0[5], N59, N156);
  xnor keyGate_0_5(N319, keyinput5, keyinput_Wire_0[5]);
  nor NOR2_34 (keyinput_Wire_0[6], N17, N42);
  xor keyGate_0_6(N322, keyinput6, keyinput_Wire_0[6]);
  and AND2_35 (keyinput_Wire_0[7], N17, N42);
  xnor keyGate_0_7(KeyNOTWire_0[3], keyinput7, keyinput_Wire_0[7]);
  not KeyNOTGate_0_3(N323, KeyNOTWire_0[3]);
nand NAND2_36 (N324, N159, N165);
or OR2_37 (N325, N159, N165);
nand NAND2_38 (N326, N171, N177);
or OR2_39 (N327, N171, N177);
nand NAND2_40 (N328, N183, N189);
or OR2_41 (N329, N183, N189);
nand NAND2_42 (N330, N195, N201);
or OR2_43 (N331, N195, N201);
and AND2_44 (N332, N210, N91);
and AND2_45 (N333, N210, N96);
and AND2_46 (N334, N210, N101);
and AND2_47 (N335, N210, N106);
and AND2_48 (N336, N210, N111);
and AND2_49 (N337, N255, N259);
and AND2_50 (N338, N210, N116);
and AND2_51 (N339, N255, N260);
and AND2_52 (N340, N210, N121);
and AND2_53 (N341, N255, N267);
not NOT1_54 (N342, N269);
not NOT1_55 (N343, N273);
or OR2_56 (N344, N270, N273);
  not NOT1_57 (keyinput_Wire_0[8], N276);
  xor keyGate_0_8(KeyNOTWire_0[4], keyinput8, keyinput_Wire_0[8]);
  not KeyNOTGate_0_4(N345, KeyNOTWire_0[4]);
not NOT1_58 (N346, N276);
  not NOT1_59 (keyinput_Wire_0[9], N279);
  xor keyGate_0_9(N347, keyinput9, keyinput_Wire_0[9]);
nor NOR2_60 (N348, N280, N284);
or OR2_61 (N349, N280, N285);
or OR2_62 (N350, N280, N286);
not NOT1_63 (N351, N293);
  not NOT1_64 (keyinput_Wire_0[10], N294);
  xor keyGate_0_10(KeyNOTWire_0[5], keyinput10, keyinput_Wire_0[10]);
  not KeyNOTGate_0_5(N352, KeyNOTWire_0[5]);
not NOT1_65 (N353, N295);
not NOT1_66 (N354, N296);
nand NAND2_67 (N355, N89, N298);
and AND2_68 (N356, N90, N298);
nand NAND2_69 (N357, N301, N302);
nand NAND2_70 (N360, N303, N304);
nand NAND2_71 (N363, N305, N306);
nand NAND2_72 (N366, N307, N308);
  not NOT1_73 (keyinput_Wire_0[11], N310);
  xor keyGate_0_11(N369, keyinput11, keyinput_Wire_0[11]);
  nor NOR2_74 (keyinput_Wire_0[12], N322, N323);
  xor keyGate_0_12(N375, keyinput12, keyinput_Wire_0[12]);
nand NAND2_75 (N376, N324, N325);
nand NAND2_76 (N379, N326, N327);
nand NAND2_77 (N382, N328, N329);
nand NAND2_78 (N385, N330, N331);
buf BUFF1_79 (N388, N290);
buf BUFF1_80 (N389, N291);
buf BUFF1_81 (N390, N292);
buf BUFF1_82 (N391, N297);
or OR2_83 (N392, N270, N343);
  not NOT1_84 (keyinput_Wire_0[13], N345);
  xnor keyGate_0_13(KeyNOTWire_0[6], keyinput13, keyinput_Wire_0[13]);
  not KeyNOTGate_0_6(N393, KeyNOTWire_0[6]);
not NOT1_85 (N399, N346);
and AND2_86 (N400, N348, N73);
not NOT1_87 (N401, N349);
not NOT1_88 (N402, N350);
not NOT1_89 (N403, N355);
not NOT1_90 (N404, N357);
not NOT1_91 (N405, N360);
and AND2_92 (N406, N357, N360);
not NOT1_93 (N407, N363);
not NOT1_94 (N408, N366);
and AND2_95 (N409, N363, N366);
  nand NAND2_96 (keyinput_Wire_0[14], N347, N352);
  xnor keyGate_0_14(N410, keyinput14, keyinput_Wire_0[14]);
not NOT1_97 (N411, N376);
not NOT1_98 (N412, N379);
and AND2_99 (N413, N376, N379);
not NOT1_100 (N414, N382);
not NOT1_101 (N415, N385);
and AND2_102 (N416, N382, N385);
and AND2_103 (N417, N210, N369);
buf BUFF1_104 (N418, N342);
buf BUFF1_105 (N419, N344);
buf BUFF1_106 (KeyWire_0_1, N351);
  xor flip_it (N420, KeyWire_0_1, KeyWire_0_2 );
buf BUFF1_107 (N421, N353);
buf BUFF1_108 (N422, N354);
buf BUFF1_109 (N423, N356);
not NOT1_110 (N424, N400);
and AND2_111 (N425, N404, N405);
and AND2_112 (N426, N407, N408);
and AND3_113 (N427, N319, N393, N55);
and AND3_114 (N432, N393, N17, N287);
  nand NAND3_115 (keyinput_Wire_0[15], N393, N287, N55);
  xor keyGate_0_15(KeyNOTWire_0[7], keyinput15, keyinput_Wire_0[15]);
  not KeyNOTGate_0_7(N437, KeyNOTWire_0[7]);
  nand NAND4_116 (keyinput_Wire_0[16], N375, N59, N156, N393);
  xnor keyGate_0_16(N442, keyinput16, keyinput_Wire_0[16]);
  nand NAND3_117 (keyinput_Wire_0[17], N393, N319, N17);
  xor keyGate_0_17(KeyNOTWire_0[8], keyinput17, keyinput_Wire_0[17]);
  not KeyNOTGate_0_8(N443, KeyNOTWire_0[8]);
and AND2_118 (N444, N411, N412);
and AND2_119 (N445, N414, N415);
buf BUFF1_120 (N446, N392);
buf BUFF1_121 (N447, N399);
buf BUFF1_122 (N448, N401);
buf BUFF1_123 (N449, N402);
buf BUFF1_124 (N450, N403);
not NOT1_125 (N451, N424);
nor NOR2_126 (N460, N406, N425);
nor NOR2_127 (N463, N409, N426);
  nand NAND2_128 (keyinput_Wire_0[18], N442, N410);
  xor keyGate_0_18(KeyNOTWire_0[9], keyinput18, keyinput_Wire_0[18]);
  not KeyNOTGate_0_9(N466, KeyNOTWire_0[9]);
and AND2_129 (N475, N143, N427);
and AND2_130 (N476, N310, N432);
and AND2_131 (N477, N146, N427);
and AND2_132 (N478, N310, N432);
and AND2_133 (N479, N149, N427);
and AND2_134 (N480, N310, N432);
and AND2_135 (N481, N153, N427);
and AND2_136 (N482, N310, N432);
  nand NAND2_137 (keyinput_Wire_0[19], N443, N1);
  xnor keyGate_0_19(N483, keyinput19, keyinput_Wire_0[19]);
or OR2_138 (N488, N369, N437);
or OR2_139 (N489, N369, N437);
or OR2_140 (N490, N369, N437);
or OR2_141 (N491, N369, N437);
nor NOR2_142 (N492, N413, N444);
nor NOR2_143 (N495, N416, N445);
nand NAND2_144 (N498, N130, N460);
or OR2_145 (N499, N130, N460);
nand NAND2_146 (N500, N463, N135);
or OR2_147 (N501, N463, N135);
and AND2_148 (N502, N91, N466);
nor NOR2_149 (N503, N475, N476);
and AND2_150 (N504, N96, N466);
nor NOR2_151 (N505, N477, N478);
and AND2_152 (N506, N101, N466);
nor NOR2_153 (N507, N479, N480);
and AND2_154 (N508, N106, N466);
nor NOR2_155 (N509, N481, N482);
and AND2_156 (N510, N143, N483);
and AND2_157 (N511, N111, N466);
and AND2_158 (N512, N146, N483);
and AND2_159 (N513, N116, N466);
and AND2_160 (N514, N149, N483);
and AND2_161 (N515, N121, N466);
and AND2_162 (N516, N153, N483);
and AND2_163 (N517, N126, N466);
nand NAND2_164 (N518, N130, N492);
or OR2_165 (N519, N130, N492);
nand NAND2_166 (N520, N495, N207);
or OR2_167 (N521, N495, N207);
and AND2_168 (N522, N451, N159);
and AND2_169 (N523, N451, N165);
and AND2_170 (N524, N451, N171);
and AND2_171 (N525, N451, N177);
and AND2_172 (N526, N451, N183);
nand NAND2_173 (N527, N451, N189);
nand NAND2_174 (N528, N451, N195);
nand NAND2_175 (N529, N451, N201);
nand NAND2_176 (N530, N498, N499);
nand NAND2_177 (N533, N500, N501);
nor NOR2_178 (N536, N309, N502);
nor NOR2_179 (N537, N316, N504);
nor NOR2_180 (N538, N317, N506);
nor NOR2_181 (N539, N318, N508);
nor NOR2_182 (N540, N510, N511);
nor NOR2_183 (N541, N512, N513);
nor NOR2_184 (N542, N514, N515);
nor NOR2_185 (N543, N516, N517);
nand NAND2_186 (N544, N518, N519);
nand NAND2_187 (N547, N520, N521);
not NOT1_188 (N550, N530);
not NOT1_189 (N551, N533);
and AND2_190 (N552, N530, N533);
nand NAND2_191 (N553, N536, N503);
nand NAND2_192 (N557, N537, N505);
nand NAND2_193 (N561, N538, N507);
nand NAND2_194 (N565, N539, N509);
nand NAND2_195 (N569, N488, N540);
nand NAND2_196 (N573, N489, N541);
nand NAND2_197 (N577, N490, N542);
  nand NAND2_198 (keyinput_Wire_0[20], N491, N543);
  xnor keyGate_0_20(N581, keyinput20, keyinput_Wire_0[20]);
not NOT1_199 (N585, N544);
not NOT1_200 (N586, N547);
and AND2_201 (N587, N544, N547);
and AND2_202 (N588, N550, N551);
and AND2_203 (N589, N585, N586);
nand NAND2_204 (N590, N553, N159);
or OR2_205 (N593, N553, N159);
and AND2_206 (N596, N246, N553);
nand NAND2_207 (N597, N557, N165);
or OR2_208 (N600, N557, N165);
and AND2_209 (N605, N246, N557);
nand NAND2_210 (N606, N561, N171);
or OR2_211 (N609, N561, N171);
and AND2_212 (N615, N246, N561);
nand NAND2_213 (N616, N565, N177);
or OR2_214 (N619, N565, N177);
and AND2_215 (N624, N246, N565);
nand NAND2_216 (N625, N569, N183);
or OR2_217 (N628, N569, N183);
and AND2_218 (N631, N246, N569);
nand NAND2_219 (N632, N573, N189);
or OR2_220 (N635, N573, N189);
and AND2_221 (N640, N246, N573);
nand NAND2_222 (N641, N577, N195);
or OR2_223 (N644, N577, N195);
and AND2_224 (N650, N246, N577);
nand NAND2_225 (N651, N581, N201);
or OR2_226 (N654, N581, N201);
and AND2_227 (N659, N246, N581);
nor NOR2_228 (N660, N552, N588);
nor NOR2_229 (N661, N587, N589);
not NOT1_230 (N662, N590);
and AND2_231 (N665, N593, N590);
nor NOR2_232 (N669, N596, N522);
not NOT1_233 (N670, N597);
and AND2_234 (N673, N600, N597);
nor NOR2_235 (N677, N605, N523);
not NOT1_236 (N678, N606);
and AND2_237 (N682, N609, N606);
nor NOR2_238 (N686, N615, N524);
not NOT1_239 (N687, N616);
and AND2_240 (N692, N619, N616);
nor NOR2_241 (N696, N624, N525);
not NOT1_242 (N697, N625);
and AND2_243 (N700, N628, N625);
nor NOR2_244 (N704, N631, N526);
not NOT1_245 (N705, N632);
and AND2_246 (N708, N635, N632);
nor NOR2_247 (N712, N337, N640);
not NOT1_248 (N713, N641);
and AND2_249 (N717, N644, N641);
nor NOR2_250 (N721, N339, N650);
not NOT1_251 (N722, N651);
and AND2_252 (N727, N654, N651);
nor NOR2_253 (N731, N341, N659);
nand NAND2_254 (N732, N654, N261);
nand NAND3_255 (N733, N644, N654, N261);
nand NAND4_256 (N734, N635, N644, N654, N261);
not NOT1_257 (N735, N662);
and AND2_258 (N736, N228, N665);
and AND2_259 (N737, N237, N662);
not NOT1_260 (N738, N670);
and AND2_261 (N739, N228, N673);
and AND2_262 (N740, N237, N670);
not NOT1_263 (N741, N678);
and AND2_264 (N742, N228, N682);
and AND2_265 (N743, N237, N678);
not NOT1_266 (N744, N687);
and AND2_267 (N745, N228, N692);
and AND2_268 (N746, N237, N687);
not NOT1_269 (N747, N697);
and AND2_270 (N748, N228, N700);
and AND2_271 (N749, N237, N697);
not NOT1_272 (N750, N705);
and AND2_273 (N751, N228, N708);
and AND2_274 (N752, N237, N705);
not NOT1_275 (N753, N713);
and AND2_276 (N754, N228, N717);
and AND2_277 (N755, N237, N713);
not NOT1_278 (N756, N722);
nor NOR2_279 (N757, N727, N261);
and AND2_280 (N758, N727, N261);
and AND2_281 (N759, N228, N727);
and AND2_282 (N760, N237, N722);
nand NAND2_283 (N761, N644, N722);
nand NAND2_284 (N762, N635, N713);
nand NAND3_285 (N763, N635, N644, N722);
nand NAND2_286 (N764, N609, N687);
nand NAND2_287 (N765, N600, N678);
nand NAND3_288 (N766, N600, N609, N687);
buf BUFF1_289 (N767, N660);
buf BUFF1_290 (N768, N661);
nor NOR2_291 (N769, N736, N737);
nor NOR2_292 (N770, N739, N740);
nor NOR2_293 (N771, N742, N743);
nor NOR2_294 (N772, N745, N746);
  nand NAND4_295 (keyinput_Wire_0[21], N750, N762, N763, N734);
  xnor keyGate_0_21(KeyNOTWire_0[10], keyinput21, keyinput_Wire_0[21]);
  not KeyNOTGate_0_10(N773, KeyNOTWire_0[10]);
nor NOR2_296 (N777, N748, N749);
nand NAND3_297 (N778, N753, N761, N733);
nor NOR2_298 (N781, N751, N752);
nand NAND2_299 (N782, N756, N732);
nor NOR2_300 (N785, N754, N755);
nor NOR2_301 (N786, N757, N758);
nor NOR2_302 (N787, N759, N760);
nor NOR2_303 (N788, N700, N773);
and AND2_304 (N789, N700, N773);
nor NOR2_305 (N790, N708, N778);
and AND2_306 (N791, N708, N778);
nor NOR2_307 (N792, N717, N782);
and AND2_308 (N793, N717, N782);
and AND2_309 (N794, N219, N786);
  nand NAND2_310 (keyinput_Wire_0[22], N628, N773);
  xnor keyGate_0_22(KeyNOTWire_0[11], keyinput22, keyinput_Wire_0[22]);
  not KeyNOTGate_0_11(N795, KeyNOTWire_0[11]);
  nand NAND2_311 (keyinput_Wire_0[23], N795, N747);
  xor keyGate_0_23(N796, keyinput23, keyinput_Wire_0[23]);
nor NOR2_312 (N802, N788, N789);
nor NOR2_313 (N803, N790, N791);
nor NOR2_314 (N804, N792, N793);
nor NOR2_315 (N805, N340, N794);
nor NOR2_316 (N806, N692, N796);
and AND2_317 (N807, N692, N796);
and AND2_318 (N808, N219, N802);
and AND2_319 (N809, N219, N803);
and AND2_320 (N810, N219, N804);
nand NAND4_321 (N811, N805, N787, N731, N529);
nand NAND2_322 (N812, N619, N796);
  nand NAND3_323 (keyinput_Wire_0[24], N609, N619, N796);
  xnor keyGate_0_24(N813, keyinput24, keyinput_Wire_0[24]);
  nand NAND4_324 (keyinput_Wire_0[25], N600, N609, N619, N796);
  xnor keyGate_0_25(KeyNOTWire_0[12], keyinput25, keyinput_Wire_0[25]);
  not KeyNOTGate_0_12(N814, KeyNOTWire_0[12]);
  nand NAND4_325 (keyinput_Wire_0[26], N738, N765, N766, N814);
  xor keyGate_0_26(KeyNOTWire_0[13], keyinput26, keyinput_Wire_0[26]);
  not KeyNOTGate_0_13(N815, KeyNOTWire_0[13]);
  nand NAND3_326 (keyinput_Wire_0[27], N741, N764, N813);
  xnor keyGate_0_27(N819, keyinput27, keyinput_Wire_0[27]);
  nand NAND2_327 (keyinput_Wire_0[28], N744, N812);
  xnor keyGate_0_28(KeyNOTWire_0[14], keyinput28, keyinput_Wire_0[28]);
  not KeyNOTGate_0_14(N822, KeyNOTWire_0[14]);
nor NOR2_328 (N825, N806, N807);
nor NOR2_329 (N826, N335, N808);
nor NOR2_330 (N827, N336, N809);
nor NOR2_331 (N828, N338, N810);
not NOT1_332 (N829, N811);
  nor NOR2_333 (keyinput_Wire_0[29], N665, N815);
  xor keyGate_0_29(KeyNOTWire_0[15], keyinput29, keyinput_Wire_0[29]);
  not KeyNOTGate_0_15(N830, KeyNOTWire_0[15]);
  and AND2_334 (keyinput_Wire_0[30], N665, N815);
  xor keyGate_0_30(KeyNOTWire_0[16], keyinput30, keyinput_Wire_0[30]);
  not KeyNOTGate_0_16(N831, KeyNOTWire_0[16]);
  nor NOR2_335 (keyinput_Wire_0[31], N673, N819);
  xnor keyGate_0_31(N832, keyinput31, keyinput_Wire_0[31]);
  and AND2_336 (keyinput_Wire_0[32], N673, N819);
  xnor keyGate_0_32(KeyNOTWire_0[17], keyinput32, keyinput_Wire_0[32]);
  not KeyNOTGate_0_17(N833, KeyNOTWire_0[17]);
  nor NOR2_337 (keyinput_Wire_0[33], N682, N822);
  xnor keyGate_0_33(N834, keyinput33, keyinput_Wire_0[33]);
  and AND2_338 (keyinput_Wire_0[34], N682, N822);
  xor keyGate_0_34(N835, keyinput34, keyinput_Wire_0[34]);
  and AND2_339 (keyinput_Wire_0[35], N219, N825);
  xnor keyGate_0_35(KeyNOTWire_0[18], keyinput35, keyinput_Wire_0[35]);
  not KeyNOTGate_0_18(N836, KeyNOTWire_0[18]);
  nand NAND3_340 (keyinput_Wire_0[36], N826, N777, N704);
  xnor keyGate_0_36(KeyNOTWire_0[19], keyinput36, keyinput_Wire_0[36]);
  not KeyNOTGate_0_19(N837, KeyNOTWire_0[19]);
nand NAND4_341 (N838, N827, N781, N712, N527);
nand NAND4_342 (N839, N828, N785, N721, N528);
not NOT1_343 (N840, N829);
  nand NAND2_344 (keyinput_Wire_0[37], N815, N593);
  xnor keyGate_0_37(KeyNOTWire_0[20], keyinput37, keyinput_Wire_0[37]);
  not KeyNOTGate_0_20(N841, KeyNOTWire_0[20]);
  nor NOR2_345 (keyinput_Wire_0[38], N830, N831);
  xor keyGate_0_38(N842, keyinput38, keyinput_Wire_0[38]);
  nor NOR2_346 (keyinput_Wire_0[39], N832, N833);
  xnor keyGate_0_39(N843, keyinput39, keyinput_Wire_0[39]);
  nor NOR2_347 (keyinput_Wire_0[40], N834, N835);
  xnor keyGate_0_40(N844, keyinput40, keyinput_Wire_0[40]);
  nor NOR2_348 (keyinput_Wire_0[41], N334, N836);
  xnor keyGate_0_41(N845, keyinput41, keyinput_Wire_0[41]);
  not NOT1_349 (keyinput_Wire_0[42], N837);
  xor keyGate_0_42(N846, keyinput42, keyinput_Wire_0[42]);
not NOT1_350 (N847, N838);
not NOT1_351 (N848, N839);
  and AND2_352 (keyinput_Wire_0[43], N735, N841);
  xor keyGate_0_43(N849, keyinput43, keyinput_Wire_0[43]);
buf BUFF1_353 (N850, N840);
  and AND2_354 (keyinput_Wire_0[44], N219, N842);
  xnor keyGate_0_44(KeyNOTWire_0[21], keyinput44, keyinput_Wire_0[44]);
  not KeyNOTGate_0_21(N851, KeyNOTWire_0[21]);
  and AND2_355 (keyinput_Wire_0[45], N219, N843);
  xnor keyGate_0_45(KeyNOTWire_0[22], keyinput45, keyinput_Wire_0[45]);
  not KeyNOTGate_0_22(N852, KeyNOTWire_0[22]);
  and AND2_356 (keyinput_Wire_0[46], N219, N844);
  xor keyGate_0_46(N853, keyinput46, keyinput_Wire_0[46]);
  nand NAND3_357 (keyinput_Wire_0[47], N845, N772, N696);
  xnor keyGate_0_47(KeyNOTWire_0[23], keyinput47, keyinput_Wire_0[47]);
  not KeyNOTGate_0_23(N854, KeyNOTWire_0[23]);
  not NOT1_358 (keyinput_Wire_0[48], N846);
  xor keyGate_0_48(KeyNOTWire_0[24], keyinput48, keyinput_Wire_0[48]);
  not KeyNOTGate_0_24(N855, KeyNOTWire_0[24]);
not NOT1_359 (N856, N847);
not NOT1_360 (N857, N848);
  not NOT1_361 (keyinput_Wire_0[49], N849);
  xor keyGate_0_49(KeyNOTWire_0[25], keyinput49, keyinput_Wire_0[49]);
  not KeyNOTGate_0_25(N858, KeyNOTWire_0[25]);
  nor NOR2_362 (keyinput_Wire_0[50], N417, N851);
  xor keyGate_0_50(N859, keyinput50, keyinput_Wire_0[50]);
  nor NOR2_363 (keyinput_Wire_0[51], N332, N852);
  xnor keyGate_0_51(N860, keyinput51, keyinput_Wire_0[51]);
  nor NOR2_364 (keyinput_Wire_0[52], N333, N853);
  xor keyGate_0_52(KeyNOTWire_0[26], keyinput52, keyinput_Wire_0[52]);
  not KeyNOTGate_0_26(N861, KeyNOTWire_0[26]);
  not NOT1_365 (keyinput_Wire_0[53], N854);
  xor keyGate_0_53(N862, keyinput53, keyinput_Wire_0[53]);
buf BUFF1_366 (N863, N855);
buf BUFF1_367 (N864, N856);
buf BUFF1_368 (N865, N857);
buf BUFF1_369 (N866, N858);
  nand NAND3_370 (keyinput_Wire_0[54], N859, N769, N669);
  xnor keyGate_0_54(N867, keyinput54, keyinput_Wire_0[54]);
  nand NAND3_371 (keyinput_Wire_0[55], N860, N770, N677);
  xor keyGate_0_55(N868, keyinput55, keyinput_Wire_0[55]);
  nand NAND3_372 (keyinput_Wire_0[56], N861, N771, N686);
  xnor keyGate_0_56(N869, keyinput56, keyinput_Wire_0[56]);
  not NOT1_373 (keyinput_Wire_0[57], N862);
  xnor keyGate_0_57(N870, keyinput57, keyinput_Wire_0[57]);
  not NOT1_374 (keyinput_Wire_0[58], N867);
  xnor keyGate_0_58(N871, keyinput58, keyinput_Wire_0[58]);
  not NOT1_375 (keyinput_Wire_0[59], N868);
  xnor keyGate_0_59(KeyNOTWire_0[27], keyinput59, keyinput_Wire_0[59]);
  not KeyNOTGate_0_27(N872, KeyNOTWire_0[27]);
  not NOT1_376 (keyinput_Wire_0[60], N869);
  xnor keyGate_0_60(N873, keyinput60, keyinput_Wire_0[60]);
buf BUFF1_377 (N874, N870);
  not NOT1_378 (keyinput_Wire_0[61], N871);
  xor keyGate_0_61(KeyNOTWire_0[28], keyinput61, keyinput_Wire_0[61]);
  not KeyNOTGate_0_28(N875, KeyNOTWire_0[28]);
  not NOT1_379 (keyinput_Wire_0[62], N872);
  xnor keyGate_0_62(N876, keyinput62, keyinput_Wire_0[62]);
  not NOT1_380 (keyinput_Wire_0[63], N873);
  xor keyGate_0_63(N877, keyinput63, keyinput_Wire_0[63]);
buf BUFF1_381 (N878, N875);
  buf BUFF1_382 (keyinput_Wire_1, N876);
  xor keyGate_1_10(N879, KeyWire_0_2, keyinput_Wire_1);
buf BUFF1_383 (N880, N877);

AntiSAT some_name( KeyWire_0_2, N207, N29, N74, N116, N138, N42, N259, N246, N96, N171, N91, N237, N126, N73, N195, N8, N101, N26, N156, N153, N159, N260, N267, N261, N177, N55, N13, N219, N89, N228, N189, N106, N1, N183, N36, N90, N201, N210, N87, N85, N80, N146, N130, N75, N86, N68, N17, N121, N255, N165, N72, N111, N135, N143, N149, N51, N152, N59, N88, N268, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183,
       keyinput184, keyinput185, keyinput186, keyinput187, keyinput188,
       keyinput189, keyinput190, keyinput191, keyinput192, keyinput193,
       keyinput194, keyinput195, keyinput196, keyinput197, keyinput198,
       keyinput199, keyinput200, keyinput201, keyinput202, keyinput203,
       keyinput204, keyinput205, keyinput206, keyinput207, keyinput208,
       keyinput209, keyinput210, keyinput211, keyinput212, keyinput213,
       keyinput214, keyinput215, keyinput216, keyinput217, keyinput218,
       keyinput219, keyinput220, keyinput221, keyinput222, keyinput223,
       keyinput224, keyinput225, keyinput226, keyinput227, keyinput228,
       keyinput229, keyinput230, keyinput231, keyinput232, keyinput233,
       keyinput234, keyinput235, keyinput236, keyinput237, keyinput238,
       keyinput239, keyinput240, keyinput241, keyinput242, keyinput243);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N207, N29, N74, N116, N138, N42, N259, N246, N96, N171, N91, N237, N126, N73, N195, N8, N101, N26, N156, N153, N159, N260, N267, N261, N177, N55, N13, N219, N89, N228, N189, N106, N1, N183, N36, N90, N201, N210, N87, N85, N80, N146, N130, N75, N86, N68, N17, N121, N255, N165, N72, N111, N135, N143, N149, N51, N152, N59, N88, N268, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183 ,
        keyinput184, keyinput185, keyinput186, keyinput187, keyinput188,
        keyinput189, keyinput190, keyinput191, keyinput192, keyinput193,
        keyinput194, keyinput195, keyinput196, keyinput197, keyinput198,
        keyinput199, keyinput200, keyinput201, keyinput202, keyinput203,
        keyinput204, keyinput205, keyinput206, keyinput207, keyinput208,
        keyinput209, keyinput210, keyinput211, keyinput212, keyinput213,
        keyinput214, keyinput215, keyinput216, keyinput217, keyinput218,
        keyinput219, keyinput220, keyinput221, keyinput222, keyinput223,
        keyinput224, keyinput225, keyinput226, keyinput227, keyinput228,
        keyinput229, keyinput230, keyinput231, keyinput232, keyinput233,
        keyinput234, keyinput235, keyinput236, keyinput237, keyinput238,
        keyinput239, keyinput240, keyinput241, keyinput242, keyinput243);

  input keyinput184, keyinput185, keyinput186, keyinput187, keyinput188;
  input keyinput189, keyinput190, keyinput191, keyinput192, keyinput193;
  input keyinput194, keyinput195, keyinput196, keyinput197, keyinput198;
  input keyinput199, keyinput200, keyinput201, keyinput202, keyinput203;
  input keyinput204, keyinput205, keyinput206, keyinput207, keyinput208;
  input keyinput209, keyinput210, keyinput211, keyinput212, keyinput213;
  input keyinput214, keyinput215, keyinput216, keyinput217, keyinput218;
  input keyinput219, keyinput220, keyinput221, keyinput222, keyinput223;
  input keyinput224, keyinput225, keyinput226, keyinput227, keyinput228;
  input keyinput229, keyinput230, keyinput231, keyinput232, keyinput233;
  input keyinput234, keyinput235, keyinput236, keyinput237, keyinput238;
  input keyinput239, keyinput240, keyinput241, keyinput242, keyinput243;

  wire [0:59] keyNTin_Wire_1;
  wire [0:28] KeyNOTWire_1;

  input N207, N29, N74, N116, N138, N42, N259, N246, N96, N171, N91, N237, N126, N73, N195, N8, N101, N26, N156, N153, N159, N260, N267, N261, N177, N55, N13, N219, N89, N228, N189, N106, N1, N183, N36, N90, N201, N210, N87, N85, N80, N146, N130, N75, N86, N68, N17, N121, N255, N165, N72, N111, N135, N143, N149, N51, N152, N59, N88, N268;
  input keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83, newWire_84, newWire_85, newWire_86, newWire_87, newWire_88, newWire_89, newWire_90, newWire_91, newWire_92, newWire_93, newWire_94, newWire_95, newWire_96, newWire_97, newWire_98, newWire_99, newWire_100, newWire_101, newWire_102, newWire_103, newWire_104, newWire_105, newWire_106, newWire_107, newWire_108, newWire_109, newWire_110, newWire_111, newWire_112, newWire_113, newWire_114, newWire_115, newWire_116, newWire_117, newWire_118, newWire_119, newWire_120, newWire_121 ;

  xnor KeyGate0 (keyNTin_Wire_1[0], N207, keyinput64);
  xor keyNTinGate_1_0(KeyNOTWire_1[0], keyinput184, keyNTin_Wire_1[0]);
  not KeyNOTGate_1_0(newWire_0, KeyNOTWire_1[0]);
  xor  KeyGate1 (newWire_1, N29, keyinput65);
  xor  KeyGate2 (newWire_2, N74, keyinput66);
  xnor KeyGate3 (newWire_3, N116, keyinput67);
  xnor KeyGate4 (keyNTin_Wire_1[1], N138, keyinput68);
  xor keyNTinGate_1_1(newWire_4, keyinput185, keyNTin_Wire_1[1]);
  xor  KeyGate5 (keyNTin_Wire_1[2], N42, keyinput69);
  xor keyNTinGate_1_2(KeyNOTWire_1[1], keyinput186, keyNTin_Wire_1[2]);
  not KeyNOTGate_1_1(newWire_5, KeyNOTWire_1[1]);
  xnor KeyGate6 (newWire_6, N259, keyinput70);
  xnor KeyGate7 (newWire_7, N246, keyinput71);
  xnor KeyGate8 (keyNTin_Wire_1[3], N96, keyinput72);
  xnor keyNTinGate_1_3(KeyNOTWire_1[2], keyinput187, keyNTin_Wire_1[3]);
  not KeyNOTGate_1_2(newWire_8, KeyNOTWire_1[2]);
  xnor KeyGate9 (newWire_9, N171, keyinput73);
  xor  KeyGate10 (keyNTin_Wire_1[4], N91, keyinput74);
  xor keyNTinGate_1_4(newWire_10, keyinput188, keyNTin_Wire_1[4]);
  xnor KeyGate11 (keyNTin_Wire_1[5], N237, keyinput75);
  xnor keyNTinGate_1_5(KeyNOTWire_1[3], keyinput189, keyNTin_Wire_1[5]);
  not KeyNOTGate_1_3(newWire_11, KeyNOTWire_1[3]);
  xor  KeyGate12 (keyNTin_Wire_1[6], N126, keyinput76);
  xor keyNTinGate_1_6(KeyNOTWire_1[4], keyinput190, keyNTin_Wire_1[6]);
  not KeyNOTGate_1_4(newWire_12, KeyNOTWire_1[4]);
  xor  KeyGate13 (newWire_13, N73, keyinput77);
  xnor KeyGate14 (keyNTin_Wire_1[7], N195, keyinput78);
  xor keyNTinGate_1_7(newWire_14, keyinput191, keyNTin_Wire_1[7]);
  xor  KeyGate15 (newWire_15, N8, keyinput79);
  xnor KeyGate16 (newWire_16, N101, keyinput80);
  xnor KeyGate17 (keyNTin_Wire_1[8], N26, keyinput81);
  xor keyNTinGate_1_8(newWire_17, keyinput192, keyNTin_Wire_1[8]);
  xnor KeyGate18 (keyNTin_Wire_1[9], N156, keyinput82);
  xor keyNTinGate_1_9(newWire_18, keyinput193, keyNTin_Wire_1[9]);
  xnor KeyGate19 (keyNTin_Wire_1[10], N153, keyinput83);
  xor keyNTinGate_1_10(KeyNOTWire_1[5], keyinput194, keyNTin_Wire_1[10]);
  not KeyNOTGate_1_5(newWire_19, KeyNOTWire_1[5]);
  xnor KeyGate20 (newWire_20, N159, keyinput84);
  xor  KeyGate21 (keyNTin_Wire_1[11], N260, keyinput85);
  xnor keyNTinGate_1_11(newWire_21, keyinput195, keyNTin_Wire_1[11]);
  xnor KeyGate22 (newWire_22, N267, keyinput86);
  xor  KeyGate23 (newWire_23, N261, keyinput87);
  xor  KeyGate24 (keyNTin_Wire_1[12], N177, keyinput88);
  xor keyNTinGate_1_12(KeyNOTWire_1[6], keyinput196, keyNTin_Wire_1[12]);
  not KeyNOTGate_1_6(newWire_24, KeyNOTWire_1[6]);
  xnor KeyGate25 (keyNTin_Wire_1[13], N55, keyinput89);
  xnor keyNTinGate_1_13(KeyNOTWire_1[7], keyinput197, keyNTin_Wire_1[13]);
  not KeyNOTGate_1_7(newWire_25, KeyNOTWire_1[7]);
  xor  KeyGate26 (keyNTin_Wire_1[14], N13, keyinput90);
  xnor keyNTinGate_1_14(KeyNOTWire_1[8], keyinput198, keyNTin_Wire_1[14]);
  not KeyNOTGate_1_8(newWire_26, KeyNOTWire_1[8]);
  xor  KeyGate27 (newWire_27, N219, keyinput91);
  xor  KeyGate28 (keyNTin_Wire_1[15], N89, keyinput92);
  xnor keyNTinGate_1_15(KeyNOTWire_1[9], keyinput199, keyNTin_Wire_1[15]);
  not KeyNOTGate_1_9(newWire_28, KeyNOTWire_1[9]);
  xnor KeyGate29 (keyNTin_Wire_1[16], N228, keyinput93);
  xnor keyNTinGate_1_16(KeyNOTWire_1[10], keyinput200, keyNTin_Wire_1[16]);
  not KeyNOTGate_1_10(newWire_29, KeyNOTWire_1[10]);
  xor  KeyGate30 (newWire_30, N189, keyinput94);
  xnor KeyGate31 (newWire_31, N106, keyinput95);
  xnor KeyGate32 (newWire_32, N1, keyinput96);
  xnor KeyGate33 (keyNTin_Wire_1[17], N183, keyinput97);
  xor keyNTinGate_1_17(newWire_33, keyinput201, keyNTin_Wire_1[17]);
  xnor KeyGate34 (newWire_34, N36, keyinput98);
  xnor KeyGate35 (keyNTin_Wire_1[18], N90, keyinput99);
  xnor keyNTinGate_1_18(newWire_35, keyinput202, keyNTin_Wire_1[18]);
  xnor KeyGate36 (newWire_36, N201, keyinput100);
  xor  KeyGate37 (newWire_37, N210, keyinput101);
  xor  KeyGate38 (newWire_38, N87, keyinput102);
  xnor KeyGate39 (keyNTin_Wire_1[19], N85, keyinput103);
  xnor keyNTinGate_1_19(KeyNOTWire_1[11], keyinput203, keyNTin_Wire_1[19]);
  not KeyNOTGate_1_11(newWire_39, KeyNOTWire_1[11]);
  xnor KeyGate40 (keyNTin_Wire_1[20], N80, keyinput104);
  xnor keyNTinGate_1_20(newWire_40, keyinput204, keyNTin_Wire_1[20]);
  xnor KeyGate41 (newWire_41, N146, keyinput105);
  xnor KeyGate42 (keyNTin_Wire_1[21], N130, keyinput106);
  xor keyNTinGate_1_21(newWire_42, keyinput205, keyNTin_Wire_1[21]);
  xor  KeyGate43 (keyNTin_Wire_1[22], N75, keyinput107);
  xor keyNTinGate_1_22(newWire_43, keyinput206, keyNTin_Wire_1[22]);
  xor  KeyGate44 (newWire_44, N86, keyinput108);
  xnor KeyGate45 (keyNTin_Wire_1[23], N68, keyinput109);
  xnor keyNTinGate_1_23(KeyNOTWire_1[12], keyinput207, keyNTin_Wire_1[23]);
  not KeyNOTGate_1_12(newWire_45, KeyNOTWire_1[12]);
  xnor KeyGate46 (newWire_46, N17, keyinput110);
  xnor KeyGate47 (keyNTin_Wire_1[24], N121, keyinput111);
  xnor keyNTinGate_1_24(newWire_47, keyinput208, keyNTin_Wire_1[24]);
  xor  KeyGate48 (newWire_48, N255, keyinput112);
  xor  KeyGate49 (newWire_49, N165, keyinput113);
  xor  KeyGate50 (newWire_50, N72, keyinput114);
  xnor KeyGate51 (newWire_51, N111, keyinput115);
  xnor KeyGate52 (newWire_52, N135, keyinput116);
  xnor KeyGate53 (keyNTin_Wire_1[25], N143, keyinput117);
  xnor keyNTinGate_1_25(newWire_53, keyinput209, keyNTin_Wire_1[25]);
  xnor KeyGate54 (keyNTin_Wire_1[26], N149, keyinput118);
  xor keyNTinGate_1_26(newWire_54, keyinput210, keyNTin_Wire_1[26]);
  xnor KeyGate55 (newWire_55, N51, keyinput119);
  xnor KeyGate56 (newWire_56, N152, keyinput120);
  xor  KeyGate57 (keyNTin_Wire_1[27], N59, keyinput121);
  xor keyNTinGate_1_27(newWire_57, keyinput211, keyNTin_Wire_1[27]);
  xor  KeyGate58 (keyNTin_Wire_1[28], N88, keyinput122);
  xor keyNTinGate_1_28(newWire_58, keyinput212, keyNTin_Wire_1[28]);
  xnor KeyGate59 (newWire_59, N268, keyinput123);
  xnor KeyGate60 (keyNTin_Wire_1[29], N207, keyinput124);
  xor keyNTinGate_1_29(newWire_60, keyinput213, keyNTin_Wire_1[29]);
  xor  KeyGate61 (keyNTin_Wire_1[30], N29, keyinput125);
  xor keyNTinGate_1_30(newWire_61, keyinput214, keyNTin_Wire_1[30]);
  xor  KeyGate62 (newWire_62, N74, keyinput126);
  xnor KeyGate63 (newWire_63, N116, keyinput127);
  xor  KeyGate64 (newWire_64, N138, keyinput128);
  xnor KeyGate65 (newWire_65, N42, keyinput129);
  xnor KeyGate66 (keyNTin_Wire_1[31], N259, keyinput130);
  xnor keyNTinGate_1_31(newWire_66, keyinput215, keyNTin_Wire_1[31]);
  xor  KeyGate67 (keyNTin_Wire_1[32], N246, keyinput131);
  xnor keyNTinGate_1_32(newWire_67, keyinput216, keyNTin_Wire_1[32]);
  xor  KeyGate68 (newWire_68, N96, keyinput132);
  xnor KeyGate69 (newWire_69, N171, keyinput133);
  xnor KeyGate70 (keyNTin_Wire_1[33], N91, keyinput134);
  xor keyNTinGate_1_33(KeyNOTWire_1[13], keyinput217, keyNTin_Wire_1[33]);
  not KeyNOTGate_1_13(newWire_70, KeyNOTWire_1[13]);
  xnor KeyGate71 (newWire_71, N237, keyinput135);
  xnor KeyGate72 (keyNTin_Wire_1[34], N126, keyinput136);
  xnor keyNTinGate_1_34(newWire_72, keyinput218, keyNTin_Wire_1[34]);
  xor  KeyGate73 (keyNTin_Wire_1[35], N73, keyinput137);
  xnor keyNTinGate_1_35(newWire_73, keyinput219, keyNTin_Wire_1[35]);
  xnor KeyGate74 (keyNTin_Wire_1[36], N195, keyinput138);
  xnor keyNTinGate_1_36(newWire_74, keyinput220, keyNTin_Wire_1[36]);
  xor  KeyGate75 (keyNTin_Wire_1[37], N8, keyinput139);
  xor keyNTinGate_1_37(newWire_75, keyinput221, keyNTin_Wire_1[37]);
  xor  KeyGate76 (newWire_76, N101, keyinput140);
  xnor KeyGate77 (newWire_77, N26, keyinput141);
  xor  KeyGate78 (newWire_78, N156, keyinput142);
  xor  KeyGate79 (newWire_79, N153, keyinput143);
  xor  KeyGate80 (newWire_80, N159, keyinput144);
  xnor KeyGate81 (keyNTin_Wire_1[38], N260, keyinput145);
  xor keyNTinGate_1_38(newWire_81, keyinput222, keyNTin_Wire_1[38]);
  xnor KeyGate82 (keyNTin_Wire_1[39], N267, keyinput146);
  xnor keyNTinGate_1_39(newWire_82, keyinput223, keyNTin_Wire_1[39]);
  xnor KeyGate83 (keyNTin_Wire_1[40], N261, keyinput147);
  xor keyNTinGate_1_40(KeyNOTWire_1[14], keyinput224, keyNTin_Wire_1[40]);
  not KeyNOTGate_1_14(newWire_83, KeyNOTWire_1[14]);
  xor  KeyGate84 (keyNTin_Wire_1[41], N177, keyinput148);
  xor keyNTinGate_1_41(newWire_84, keyinput225, keyNTin_Wire_1[41]);
  xnor KeyGate85 (newWire_85, N55, keyinput149);
  xnor KeyGate86 (newWire_86, N13, keyinput150);
  xor  KeyGate87 (newWire_87, N219, keyinput151);
  xnor KeyGate88 (keyNTin_Wire_1[42], N89, keyinput152);
  xor keyNTinGate_1_42(newWire_88, keyinput226, keyNTin_Wire_1[42]);
  xor  KeyGate89 (keyNTin_Wire_1[43], N228, keyinput153);
  xor keyNTinGate_1_43(KeyNOTWire_1[15], keyinput227, keyNTin_Wire_1[43]);
  not KeyNOTGate_1_15(newWire_89, KeyNOTWire_1[15]);
  xnor KeyGate90 (keyNTin_Wire_1[44], N189, keyinput154);
  xnor keyNTinGate_1_44(newWire_90, keyinput228, keyNTin_Wire_1[44]);
  xor  KeyGate91 (keyNTin_Wire_1[45], N106, keyinput155);
  xnor keyNTinGate_1_45(KeyNOTWire_1[16], keyinput229, keyNTin_Wire_1[45]);
  not KeyNOTGate_1_16(newWire_91, KeyNOTWire_1[16]);
  xor  KeyGate92 (newWire_92, N1, keyinput156);
  xor  KeyGate93 (keyNTin_Wire_1[46], N183, keyinput157);
  xnor keyNTinGate_1_46(newWire_93, keyinput230, keyNTin_Wire_1[46]);
  xnor KeyGate94 (keyNTin_Wire_1[47], N36, keyinput158);
  xor keyNTinGate_1_47(KeyNOTWire_1[17], keyinput231, keyNTin_Wire_1[47]);
  not KeyNOTGate_1_17(newWire_94, KeyNOTWire_1[17]);
  xnor KeyGate95 (keyNTin_Wire_1[48], N90, keyinput159);
  xnor keyNTinGate_1_48(KeyNOTWire_1[18], keyinput232, keyNTin_Wire_1[48]);
  not KeyNOTGate_1_18(newWire_95, KeyNOTWire_1[18]);
  xor  KeyGate96 (newWire_96, N201, keyinput160);
  xnor KeyGate97 (newWire_97, N210, keyinput161);
  xnor KeyGate98 (newWire_98, N87, keyinput162);
  xor  KeyGate99 (newWire_99, N85, keyinput163);
  xnor KeyGate100 (newWire_100, N80, keyinput164);
  xor  KeyGate101 (newWire_101, N146, keyinput165);
  xor  KeyGate102 (newWire_102, N130, keyinput166);
  xor  KeyGate103 (keyNTin_Wire_1[49], N75, keyinput167);
  xnor keyNTinGate_1_49(KeyNOTWire_1[19], keyinput233, keyNTin_Wire_1[49]);
  not KeyNOTGate_1_19(newWire_103, KeyNOTWire_1[19]);
  xor  KeyGate104 (keyNTin_Wire_1[50], N86, keyinput168);
  xor keyNTinGate_1_50(newWire_104, keyinput234, keyNTin_Wire_1[50]);
  xor  KeyGate105 (keyNTin_Wire_1[51], N68, keyinput169);
  xnor keyNTinGate_1_51(KeyNOTWire_1[20], keyinput235, keyNTin_Wire_1[51]);
  not KeyNOTGate_1_20(newWire_105, KeyNOTWire_1[20]);
  xor  KeyGate106 (newWire_106, N17, keyinput170);
  xnor KeyGate107 (keyNTin_Wire_1[52], N121, keyinput171);
  xor keyNTinGate_1_52(KeyNOTWire_1[21], keyinput236, keyNTin_Wire_1[52]);
  not KeyNOTGate_1_21(newWire_107, KeyNOTWire_1[21]);
  xor  KeyGate108 (newWire_108, N255, keyinput172);
  xnor KeyGate109 (newWire_109, N165, keyinput173);
  xor  KeyGate110 (newWire_110, N72, keyinput174);
  xnor KeyGate111 (newWire_111, N111, keyinput175);
  xor  KeyGate112 (newWire_112, N135, keyinput176);
  xor  KeyGate113 (keyNTin_Wire_1[53], N143, keyinput177);
  xor keyNTinGate_1_53(KeyNOTWire_1[22], keyinput237, keyNTin_Wire_1[53]);
  not KeyNOTGate_1_22(newWire_113, KeyNOTWire_1[22]);
  xor  KeyGate114 (newWire_114, N149, keyinput178);
  xnor KeyGate115 (keyNTin_Wire_1[54], N51, keyinput179);
  xor keyNTinGate_1_54(KeyNOTWire_1[23], keyinput238, keyNTin_Wire_1[54]);
  not KeyNOTGate_1_23(newWire_115, KeyNOTWire_1[23]);
  xnor KeyGate116 (keyNTin_Wire_1[55], N152, keyinput180);
  xnor keyNTinGate_1_55(KeyNOTWire_1[24], keyinput239, keyNTin_Wire_1[55]);
  not KeyNOTGate_1_24(newWire_116, KeyNOTWire_1[24]);
  xor  KeyGate117 (keyNTin_Wire_1[56], N59, keyinput181);
  xor keyNTinGate_1_56(KeyNOTWire_1[25], keyinput240, keyNTin_Wire_1[56]);
  not KeyNOTGate_1_25(newWire_117, KeyNOTWire_1[25]);
  xor  KeyGate118 (keyNTin_Wire_1[57], N88, keyinput182);
  xor keyNTinGate_1_57(KeyNOTWire_1[26], keyinput241, keyNTin_Wire_1[57]);
  not KeyNOTGate_1_26(newWire_118, KeyNOTWire_1[26]);
  xor  KeyGate119 (keyNTin_Wire_1[58], N268, keyinput183);
  xor keyNTinGate_1_58(KeyNOTWire_1[27], keyinput242, keyNTin_Wire_1[58]);
  not KeyNOTGate_1_27(newWire_119, KeyNOTWire_1[27]);
  and some_function (newWire_120, newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59 );
  nand compl_function (keyNTin_Wire_1[59], newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83, newWire_84, newWire_85, newWire_86, newWire_87, newWire_88, newWire_89, newWire_90, newWire_91, newWire_92, newWire_93, newWire_94, newWire_95, newWire_96, newWire_97, newWire_98, newWire_99, newWire_100, newWire_101, newWire_102, newWire_103, newWire_104, newWire_105, newWire_106, newWire_107, newWire_108, newWire_109, newWire_110, newWire_111, newWire_112, newWire_113, newWire_114, newWire_115, newWire_116, newWire_117, newWire_118, newWire_119);
  xor keyNTinGate_1_59(KeyNOTWire_1[28], keyinput243, keyNTin_Wire_1[59]);
  not KeyNOTGate_1_28(newWire_121, KeyNOTWire_1[28]);
  and finalAND (KeyWire_0_2, newWire_120, newWire_121);

endmodule /* AntiSAT */
