// Verilog File 
module top (G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,
G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,
G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,
G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat,G223gat,G329gat,G370gat,
G421gat,G430gat,G431gat,G432gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,
keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,
keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,
keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,keyinput35,
keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,keyinput45,
keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52);

input G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,
G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,
G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,
G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat,keyinput0,keyinput1,keyinput2,
keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,
keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,
keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,
keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,
keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52;

output G223gat,G329gat,G370gat,G421gat,G430gat,G431gat,G432gat;

wire G118gat,G119gat,G122gat,G123gat,G126gat,G127gat,G130gat,G131gat,G134gat,
G135gat,G138gat,G139gat,G142gat,G143gat,G146gat,G147gat,G150gat,G151gat,G154gat,
G157gat,G158gat,G159gat,G162gat,G165gat,G168gat,G171gat,G174gat,G177gat,G180gat,
G183gat,G184gat,G185gat,G186gat,G187gat,G188gat,G189gat,G190gat,G191gat,G192gat,
G193gat,G194gat,G195gat,G196gat,G197gat,G198gat,G199gat,G203gat,G213gat,G224gat,
G227gat,G230gat,G233gat,G236gat,G239gat,G242gat,G243gat,G246gat,G247gat,G250gat,
G251gat,G254gat,G255gat,G256gat,G257gat,G258gat,G259gat,G260gat,G263gat,G264gat,
G267gat,G270gat,G273gat,G276gat,G279gat,G282gat,G285gat,G288gat,G289gat,G290gat,
G291gat,G292gat,G293gat,G294gat,G295gat,G296gat,G300gat,G301gat,G302gat,G303gat,
G304gat,G305gat,G306gat,G307gat,G308gat,G309gat,G319gat,G330gat,G331gat,G332gat,
G333gat,G334gat,G335gat,G336gat,G337gat,G338gat,G339gat,G340gat,G341gat,G342gat,
G343gat,G344gat,G345gat,G346gat,G347gat,G348gat,G349gat,G350gat,G351gat,G352gat,
G353gat,G354gat,G355gat,G356gat,G357gat,G360gat,G371gat,G372gat,G373gat,G374gat,
G375gat,G376gat,G377gat,G378gat,G379gat,G380gat,G381gat,G386gat,G393gat,G399gat,
G404gat,G407gat,G411gat,G414gat,G415gat,G416gat,G417gat,G418gat,G419gat,G420gat,
G422gat,G425gat,G428gat,G429gat,muxed0,muxed1,muxed2,muxed3,muxed4,muxed5,
muxed6,muxed7,muxed8,muxed9,muxed10,muxed11,muxed12,muxed13,muxed14,muxed15,
muxed16,muxed17,muxed18,muxed19,muxed20,muxed21,muxed22,muxed23,muxed24,muxed25,
muxed26,muxed27,muxed28,muxed29,muxed30,muxed31,muxed32,muxed33,muxed34,muxed35,
muxed36,muxed37,muxed38,muxed39,muxed40,muxed41,muxed42,muxed43,muxed44,muxed45,
muxed46,muxed47,muxed48,muxed49,muxed50,muxed51,muxed52;
not gate_0(G118gat,G1gat);
not gate_1(G119gat,G4gat);
not gate_2(G122gat,G11gat);
not gate_3(G123gat,G17gat);
not gate_4(G126gat,G24gat);
not gate_5(G127gat,G30gat);
not gate_6(G130gat,G37gat);
not gate_7(G131gat,G43gat);
not gate_8(G134gat,G50gat);
not gate_9(G135gat,G56gat);
not gate_10(G138gat,G63gat);
not gate_11(G139gat,G69gat);
not gate_12(G142gat,G76gat);
not gate_13(G143gat,G82gat);
not gate_14(G146gat,G89gat);
not gate_15(G147gat,G95gat);
not gate_16(G150gat,G102gat);
not gate_17(G151gat,G108gat);
nand gate_18(G154gat,G118gat,G4gat);
nor gate_19(G157gat,G8gat,G119gat);
nor gate_20(G158gat,G14gat,G119gat);
nand gate_21(G159gat,muxed43,G17gat);
nand gate_22(G162gat,G126gat,G30gat);
nand gate_23(G165gat,G130gat,G43gat);
nand gate_24(G168gat,G134gat,G56gat);
nand gate_25(G171gat,G138gat,G69gat);
nand gate_26(G174gat,muxed21,G82gat);
nand gate_27(G177gat,G146gat,G95gat);
nand gate_28(G180gat,G150gat,G108gat);
nor gate_29(G183gat,G21gat,G123gat);
nor gate_30(G184gat,G27gat,G123gat);
nor gate_31(G185gat,G34gat,G127gat);
nor gate_32(G186gat,G40gat,G127gat);
nor gate_33(G187gat,G47gat,G131gat);
nor gate_34(G188gat,G53gat,G131gat);
nor gate_35(G189gat,G60gat,G135gat);
nor gate_36(G190gat,G66gat,G135gat);
nor gate_37(G191gat,G73gat,G139gat);
nor gate_38(G192gat,G79gat,G139gat);
nor gate_39(G193gat,G86gat,G143gat);
nor gate_40(G194gat,G92gat,G143gat);
nor gate_41(G195gat,G99gat,G147gat);
nor gate_42(G196gat,G105gat,G147gat);
nor gate_43(G197gat,G112gat,G151gat);
nor gate_44(G198gat,G115gat,G151gat);
and gate_45(G199gat,G154gat,muxed42,G162gat,G165gat,G168gat,G171gat,G174gat,G177gat,G180gat);
not gate_46(G203gat,G199gat);
not gate_47(G213gat,G199gat);
not gate_48(G223gat,G199gat);
xor gate_49(G224gat,G203gat,G154gat);
xor gate_50(G227gat,G203gat,muxed42);
xor gate_51(G230gat,G203gat,G162gat);
xor gate_52(G233gat,G203gat,G165gat);
xor gate_53(G236gat,G203gat,G168gat);
xor gate_54(G239gat,G203gat,G171gat);
nand gate_55(G242gat,G1gat,muxed48);
xor gate_56(G243gat,G203gat,G174gat);
nand gate_57(G246gat,muxed48,G11gat);
xor gate_58(G247gat,G203gat,G177gat);
nand gate_59(G250gat,muxed48,G24gat);
xor gate_60(G251gat,G203gat,G180gat);
nand gate_61(G254gat,muxed48,G37gat);
nand gate_62(G255gat,muxed48,G50gat);
nand gate_63(G256gat,muxed48,G63gat);
nand gate_64(G257gat,muxed48,G76gat);
nand gate_65(G258gat,muxed48,G89gat);
nand gate_66(G259gat,muxed48,G102gat);
nand gate_67(G260gat,G224gat,muxed25);
nand gate_68(G263gat,G224gat,G158gat);
nand gate_69(G264gat,muxed41,G183gat);
nand gate_70(G267gat,G230gat,muxed50);
nand gate_71(G270gat,G233gat,muxed23);
nand gate_72(G273gat,G236gat,G189gat);
nand gate_73(G276gat,G239gat,G191gat);
nand gate_74(G279gat,G243gat,G193gat);
nand gate_75(G282gat,G247gat,muxed9);
nand gate_76(G285gat,G251gat,G197gat);
nand gate_77(G288gat,muxed41,G184gat);
nand gate_78(G289gat,G230gat,muxed33);
nand gate_79(G290gat,G233gat,G188gat);
nand gate_80(G291gat,G236gat,G190gat);
nand gate_81(G292gat,G239gat,G192gat);
nand gate_82(G293gat,G243gat,G194gat);
nand gate_83(G294gat,G247gat,G196gat);
nand gate_84(G295gat,G251gat,muxed4);
and gate_85(G296gat,muxed24,G264gat,G267gat,G270gat,G273gat,G276gat,G279gat,G282gat,G285gat);
not gate_86(G300gat,G263gat);
not gate_87(G301gat,G288gat);
not gate_88(G302gat,G289gat);
not gate_89(G303gat,G290gat);
not gate_90(G304gat,G291gat);
not gate_91(G305gat,G292gat);
not gate_92(G306gat,G293gat);
not gate_93(G307gat,muxed40);
not gate_94(G308gat,muxed39);
not gate_95(G309gat,muxed2);
not gate_96(G319gat,muxed2);
not gate_97(G329gat,muxed2);
xor gate_98(G330gat,muxed28,muxed24);
xor gate_99(G331gat,muxed28,G264gat);
xor gate_100(G332gat,muxed28,G267gat);
xor gate_101(G333gat,muxed28,G270gat);
nand gate_102(G334gat,G8gat,G319gat);
xor gate_103(G335gat,muxed28,G273gat);
nand gate_104(G336gat,G319gat,G21gat);
xor gate_105(G337gat,muxed28,G276gat);
nand gate_106(G338gat,G319gat,G34gat);
xor gate_107(G339gat,muxed28,G279gat);
nand gate_108(G340gat,G319gat,G47gat);
xor gate_109(G341gat,muxed28,G282gat);
nand gate_110(G342gat,G319gat,G60gat);
xor gate_111(G343gat,muxed28,G285gat);
nand gate_112(G344gat,G319gat,G73gat);
nand gate_113(G345gat,G319gat,G86gat);
nand gate_114(G346gat,G319gat,G99gat);
nand gate_115(G347gat,G319gat,G112gat);
nand gate_116(G348gat,muxed52,G300gat);
nand gate_117(G349gat,G331gat,G301gat);
nand gate_118(G350gat,G332gat,G302gat);
nand gate_119(G351gat,muxed38,G303gat);
nand gate_120(G352gat,muxed0,G304gat);
nand gate_121(G353gat,muxed44,G305gat);
nand gate_122(G354gat,G339gat,G306gat);
nand gate_123(G355gat,G341gat,muxed51);
nand gate_124(G356gat,muxed19,G308gat);
and gate_125(G357gat,muxed20,G349gat,G350gat,muxed37,muxed12,G353gat,muxed13,muxed49,G356gat);
not gate_126(G360gat,muxed31);
not gate_127(G370gat,muxed31);
nand gate_128(G371gat,G14gat,muxed10);
nand gate_129(G372gat,muxed10,G27gat);
nand gate_130(G373gat,muxed10,G40gat);
nand gate_131(G374gat,muxed10,G53gat);
nand gate_132(G375gat,muxed10,G66gat);
nand gate_133(G376gat,muxed10,G79gat);
nand gate_134(G377gat,muxed10,G92gat);
nand gate_135(G378gat,muxed10,G105gat);
nand gate_136(G379gat,muxed10,G115gat);
nand gate_137(G380gat,G4gat,G242gat,G334gat,G371gat);
nand gate_138(G381gat,G246gat,G336gat,G372gat,G17gat);
nand gate_139(G386gat,muxed29,G338gat,G373gat,G30gat);
nand gate_140(G393gat,G254gat,G340gat,G374gat,G43gat);
nand gate_141(G399gat,G255gat,G342gat,G375gat,G56gat);
nand gate_142(G404gat,G256gat,G344gat,G376gat,G69gat);
nand gate_143(G407gat,G257gat,G345gat,G377gat,G82gat);
nand gate_144(G411gat,G258gat,G346gat,muxed8,G95gat);
nand gate_145(G414gat,G259gat,G347gat,G379gat,G108gat);
not gate_146(G415gat,G380gat);
and gate_147(G416gat,G381gat,G386gat,G393gat,G399gat,G404gat,G407gat,muxed14,G414gat);
not gate_148(G417gat,G393gat);
not gate_149(G418gat,G404gat);
not gate_150(G419gat,G407gat);
not gate_151(G420gat,muxed14);
nor gate_152(G421gat,G415gat,G416gat);
nand gate_153(G422gat,G386gat,G417gat);
nand gate_154(G425gat,G386gat,G393gat,G418gat,G399gat);
nand gate_155(G428gat,G399gat,G393gat,G419gat);
nand gate_156(G429gat,G386gat,G393gat,G407gat,muxed5);
nand gate_157(G430gat,G381gat,G386gat,G422gat,G399gat);
nand gate_158(G431gat,G381gat,G386gat,G425gat,G428gat);
nand gate_159(G432gat,G381gat,G422gat,G425gat,muxed3);
assign muxed0 = keyinput0 ? G335gat : muxed1;
assign muxed1 = keyinput1 ? G432gat : G184gat;
assign muxed2 = keyinput2 ? G296gat : G432gat;
assign muxed3 = keyinput3 ? G429gat : G296gat;
assign muxed4 = keyinput4 ? G198gat : G429gat;
assign muxed5 = keyinput5 ? muxed27 : G224gat;
assign muxed6 = keyinput6 ? G157gat : muxed27;
assign muxed7 = keyinput7 ? G411gat : G371gat;
assign muxed8 = keyinput8 ? G378gat : G191gat;
assign muxed9 = keyinput9 ? G195gat : G378gat;
assign muxed10 = keyinput10 ? G360gat : G338gat;
assign muxed11 = keyinput11 ? muxed34 : G192gat;
assign muxed12 = keyinput12 ? G352gat : muxed37;
assign muxed13 = keyinput13 ? G354gat : G352gat;
assign muxed14 = keyinput14 ? muxed7 : muxed15;
assign muxed15 = keyinput15 ? muxed30 : G171gat;
assign muxed16 = keyinput16 ? G250gat : muxed30;
assign muxed17 = keyinput17 ? muxed32 : G422gat;
assign muxed18 = keyinput18 ? muxed46 : G360gat;
assign muxed19 = keyinput19 ? G343gat : muxed46;
assign muxed20 = keyinput20 ? G348gat : G304gat;
assign muxed21 = keyinput21 ? G142gat : G348gat;
assign muxed22 = keyinput22 ? G330gat : G190gat;
assign muxed23 = keyinput23 ? G187gat : G330gat;
assign muxed24 = keyinput24 ? G260gat : G296gat;
assign muxed25 = keyinput25 ? muxed26 : G302gat;
assign muxed26 = keyinput26 ? muxed6 : muxed6;
assign muxed27 = keyinput27 ? G420gat : G296gat;
assign muxed28 = keyinput28 ? G309gat : muxed29;
assign muxed29 = keyinput29 ? muxed16 : muxed40;
assign muxed30 = keyinput30 ? G370gat : G422gat;
assign muxed31 = keyinput31 ? muxed17 : G126gat;
assign muxed32 = keyinput32 ? muxed11 : muxed37;
assign muxed33 = keyinput33 ? G186gat : muxed11;
assign muxed34 = keyinput34 ? muxed45 : muxed42;
assign muxed35 = keyinput35 ? G122gat : muxed45;
assign muxed36 = keyinput36 ? muxed47 : G239gat;
assign muxed37 = keyinput37 ? G351gat : muxed7;
assign muxed38 = keyinput38 ? G333gat : G353gat;
assign muxed39 = keyinput39 ? G295gat : G333gat;
assign muxed40 = keyinput40 ? G294gat : muxed41;
assign muxed41 = keyinput41 ? G227gat : G399gat;
assign muxed42 = keyinput42 ? G159gat : G282gat;
assign muxed43 = keyinput43 ? muxed35 : G270gat;
assign muxed44 = keyinput44 ? G337gat : muxed35;
assign muxed45 = keyinput45 ? muxed18 : G319gat;
assign muxed46 = keyinput46 ? muxed36 : muxed14;
assign muxed47 = keyinput47 ? G357gat : G247gat;
assign muxed48 = keyinput48 ? G213gat : G357gat;
assign muxed49 = keyinput49 ? G355gat : G146gat;
assign muxed50 = keyinput50 ? G185gat : G355gat;
assign muxed51 = keyinput51 ? G307gat : G138gat;
assign muxed52 = keyinput52 ? muxed22 : G307gat;
endmodule
