`timescale 1ns / 1ps
// Verilog
// c432
// Ninputs 36
// Noutputs 7
// NtotalGates 160
// NOT1 40
// NAND2 64
// NOR2 19
// AND9 3
// XOR2 18
// NAND4 14
// AND8 1
// NAND3 1

module top (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
                  N430,N431,N432,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
                  keyinput30, keyinput31,
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36,
        keyinput37, keyinput38, keyinput39, keyinput40, keyinput41,
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46,
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51,
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56,
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61,
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66,
        keyinput67, keyinput68, keyinput69, keyinput70, keyinput71,
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76,
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81,
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86,
        keyinput87, keyinput88, keyinput89, keyinput90, keyinput91,
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96,
        keyinput97, keyinput98, keyinput99, keyinput100, keyinput101,
                  keyinput102, keyinput103,
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
        keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
        keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
        keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
        keyinput139);

  input keyinput104, keyinput105, keyinput106, keyinput107, keyinput108;
  input keyinput109, keyinput110, keyinput111, keyinput112, keyinput113;
  input keyinput114, keyinput115, keyinput116, keyinput117, keyinput118;
  input keyinput119, keyinput120, keyinput121, keyinput122, keyinput123;
  input keyinput124, keyinput125, keyinput126, keyinput127, keyinput128;
  input keyinput129, keyinput130, keyinput131, keyinput132, keyinput133;
  input keyinput134, keyinput135, keyinput136, keyinput137, keyinput138;
  input keyinput139;


  input keyinput32, keyinput33, keyinput34, keyinput35, keyinput36;
  input keyinput37, keyinput38, keyinput39, keyinput40, keyinput41;
  input keyinput42, keyinput43, keyinput44, keyinput45, keyinput46;
  input keyinput47, keyinput48, keyinput49, keyinput50, keyinput51;
  input keyinput52, keyinput53, keyinput54, keyinput55, keyinput56;
  input keyinput57, keyinput58, keyinput59, keyinput60, keyinput61;
  input keyinput62, keyinput63, keyinput64, keyinput65, keyinput66;
  input keyinput67, keyinput68, keyinput69, keyinput70, keyinput71;
  input keyinput72, keyinput73, keyinput74, keyinput75, keyinput76;
  input keyinput77, keyinput78, keyinput79, keyinput80, keyinput81;
  input keyinput82, keyinput83, keyinput84, keyinput85, keyinput86;
  input keyinput87, keyinput88, keyinput89, keyinput90, keyinput91;
  input keyinput92, keyinput93, keyinput94, keyinput95, keyinput96;
  input keyinput97, keyinput98, keyinput99, keyinput100, keyinput101;
  input keyinput102, keyinput103;

  wire KeyWire_0_1 , KeyWire_0_2;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31;

  wire [0:31] keyinput_Wire_0;
  wire [0:17] KeyNOTWire_0;

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;

output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429;

  not NOT1_1 (keyinput_Wire_0[0], N1);
  xnor keyGate_0_0(N118, keyinput0, keyinput_Wire_0[0]);
not NOT1_2 (N119, N4);
  not NOT1_3 (keyinput_Wire_0[1], N11);
  xnor keyGate_0_1(N122, keyinput1, keyinput_Wire_0[1]);
not NOT1_4 (N123, N17);
  not NOT1_5 (keyinput_Wire_0[2], N24);
  xor keyGate_0_2(N126, keyinput2, keyinput_Wire_0[2]);
not NOT1_6 (N127, N30);
  not NOT1_7 (keyinput_Wire_0[3], N37);
  xnor keyGate_0_3(KeyNOTWire_0[0], keyinput3, keyinput_Wire_0[3]);
  not KeyNOTGate_0_0(N130, KeyNOTWire_0[0]);
not NOT1_8 (N131, N43);
  not NOT1_9 (keyinput_Wire_0[4], N50);
  xor keyGate_0_4(KeyNOTWire_0[1], keyinput4, keyinput_Wire_0[4]);
  not KeyNOTGate_0_1(N134, KeyNOTWire_0[1]);
not NOT1_10 (N135, N56);
  not NOT1_11 (keyinput_Wire_0[5], N63);
  xor keyGate_0_5(N138, keyinput5, keyinput_Wire_0[5]);
not NOT1_12 (N139, N69);
  not NOT1_13 (keyinput_Wire_0[6], N76);
  xnor keyGate_0_6(N142, keyinput6, keyinput_Wire_0[6]);
not NOT1_14 (N143, N82);
  not NOT1_15 (keyinput_Wire_0[7], N89);
  xor keyGate_0_7(N146, keyinput7, keyinput_Wire_0[7]);
not NOT1_16 (N147, N95);
  not NOT1_17 (keyinput_Wire_0[8], N102);
  xnor keyGate_0_8(KeyNOTWire_0[2], keyinput8, keyinput_Wire_0[8]);
  not KeyNOTGate_0_2(N150, KeyNOTWire_0[2]);
not NOT1_18 (N151, N108);
  nand NAND2_19 (keyinput_Wire_0[9], N118, N4);
  xnor keyGate_0_9(KeyNOTWire_0[3], keyinput9, keyinput_Wire_0[9]);
  not KeyNOTGate_0_3(N154, KeyNOTWire_0[3]);
nor NOR2_20 (N157, N8, N119);
nor NOR2_21 (N158, N14, N119);
  nand NAND2_22 (keyinput_Wire_0[10], N122, N17);
  xnor keyGate_0_10(KeyNOTWire_0[4], keyinput10, keyinput_Wire_0[10]);
  not KeyNOTGate_0_4(N159, KeyNOTWire_0[4]);
  nand NAND2_23 (keyinput_Wire_0[11], N126, N30);
  xnor keyGate_0_11(KeyNOTWire_0[5], keyinput11, keyinput_Wire_0[11]);
  not KeyNOTGate_0_5(N162, KeyNOTWire_0[5]);
  nand NAND2_24 (keyinput_Wire_0[12], N130, N43);
  xnor keyGate_0_12(N165, keyinput12, keyinput_Wire_0[12]);
  nand NAND2_25 (keyinput_Wire_0[13], N134, N56);
  xnor keyGate_0_13(KeyNOTWire_0[6], keyinput13, keyinput_Wire_0[13]);
  not KeyNOTGate_0_6(N168, KeyNOTWire_0[6]);
  nand NAND2_26 (keyinput_Wire_0[14], N138, N69);
  xnor keyGate_0_14(KeyNOTWire_0[7], keyinput14, keyinput_Wire_0[14]);
  not KeyNOTGate_0_7(N171, KeyNOTWire_0[7]);
  nand NAND2_27 (keyinput_Wire_0[15], N142, N82);
  xnor keyGate_0_15(KeyNOTWire_0[8], keyinput15, keyinput_Wire_0[15]);
  not KeyNOTGate_0_8(N174, KeyNOTWire_0[8]);
  nand NAND2_28 (keyinput_Wire_0[16], N146, N95);
  xor keyGate_0_16(KeyNOTWire_0[9], keyinput16, keyinput_Wire_0[16]);
  not KeyNOTGate_0_9(N177, KeyNOTWire_0[9]);
  nand NAND2_29 (keyinput_Wire_0[17], N150, N108);
  xnor keyGate_0_17(KeyNOTWire_0[10], keyinput17, keyinput_Wire_0[17]);
  not KeyNOTGate_0_10(N180, KeyNOTWire_0[10]);
nor NOR2_30 (N183, N21, N123);
nor NOR2_31 (N184, N27, N123);
nor NOR2_32 (N185, N34, N127);
nor NOR2_33 (N186, N40, N127);
nor NOR2_34 (N187, N47, N131);
nor NOR2_35 (N188, N53, N131);
nor NOR2_36 (N189, N60, N135);
nor NOR2_37 (N190, N66, N135);
nor NOR2_38 (N191, N73, N139);
nor NOR2_39 (N192, N79, N139);
nor NOR2_40 (N193, N86, N143);
nor NOR2_41 (N194, N92, N143);
nor NOR2_42 (N195, N99, N147);
nor NOR2_43 (N196, N105, N147);
nor NOR2_44 (N197, N112, N151);
nor NOR2_45 (N198, N115, N151);
  and AND9_46 (keyinput_Wire_0[18], N154, N159, N162, N165, N168, N171, N174, N177, N180);
  xnor keyGate_0_18(KeyNOTWire_0[11], keyinput18, keyinput_Wire_0[18]);
  not KeyNOTGate_0_11(N199, KeyNOTWire_0[11]);
  not NOT1_47 (keyinput_Wire_0[19], N199);
  xnor keyGate_0_19(N203, keyinput19, keyinput_Wire_0[19]);
not NOT1_48 (N213, N199);
not NOT1_49 (N223, N199);
xor XOR2_50 (N224, N203, N154);
xor XOR2_51 (N227, N203, N159);
xor XOR2_52 (N230, N203, N162);
xor XOR2_53 (N233, N203, N165);
xor XOR2_54 (N236, N203, N168);
xor XOR2_55 (N239, N203, N171);
nand NAND2_56 (N242, N1, N213);
xor XOR2_57 (N243, N203, N174);
nand NAND2_58 (N246, N213, N11);
xor XOR2_59 (N247, N203, N177);
nand NAND2_60 (N250, N213, N24);
xor XOR2_61 (N251, N203, N180);
nand NAND2_62 (N254, N213, N37);
nand NAND2_63 (N255, N213, N50);
nand NAND2_64 (N256, N213, N63);
nand NAND2_65 (N257, N213, N76);
nand NAND2_66 (N258, N213, N89);
nand NAND2_67 (N259, N213, N102);
nand NAND2_68 (N260, N224, N157);
nand NAND2_69 (N263, N224, N158);
nand NAND2_70 (N264, N227, N183);
nand NAND2_71 (N267, N230, N185);
nand NAND2_72 (N270, N233, N187);
nand NAND2_73 (N273, N236, N189);
nand NAND2_74 (N276, N239, N191);
nand NAND2_75 (N279, N243, N193);
nand NAND2_76 (N282, N247, N195);
nand NAND2_77 (N285, N251, N197);
nand NAND2_78 (N288, N227, N184);
nand NAND2_79 (N289, N230, N186);
nand NAND2_80 (N290, N233, N188);
nand NAND2_81 (N291, N236, N190);
nand NAND2_82 (N292, N239, N192);
nand NAND2_83 (N293, N243, N194);
nand NAND2_84 (N294, N247, N196);
nand NAND2_85 (N295, N251, N198);
  and AND9_86 (keyinput_Wire_0[20], N260, N264, N267, N270, N273, N276, N279, N282, N285);
  xor keyGate_0_20(N296, keyinput20, keyinput_Wire_0[20]);
not NOT1_87 (N300, N263);
not NOT1_88 (N301, N288);
not NOT1_89 (N302, N289);
not NOT1_90 (N303, N290);
not NOT1_91 (N304, N291);
not NOT1_92 (N305, N292);
not NOT1_93 (N306, N293);
not NOT1_94 (N307, N294);
not NOT1_95 (N308, N295);
  not NOT1_96 (keyinput_Wire_0[21], N296);
  xor keyGate_0_21(KeyNOTWire_0[12], keyinput21, keyinput_Wire_0[21]);
  not KeyNOTGate_0_12(N309, KeyNOTWire_0[12]);
not NOT1_97 (N319, N296);
not NOT1_98 (N329, N296);
xor XOR2_99 (N330, N309, N260);
xor XOR2_100 (N331, N309, N264);
xor XOR2_101 (N332, N309, N267);
xor XOR2_102 (N333, N309, N270);
nand NAND2_103 (N334, N8, N319);
xor XOR2_104 (N335, N309, N273);
nand NAND2_105 (N336, N319, N21);
xor XOR2_106 (N337, N309, N276);
nand NAND2_107 (N338, N319, N34);
xor XOR2_108 (N339, N309, N279);
nand NAND2_109 (N340, N319, N47);
xor XOR2_110 (N341, N309, N282);
nand NAND2_111 (N342, N319, N60);
xor XOR2_112 (N343, N309, N285);
nand NAND2_113 (N344, N319, N73);
nand NAND2_114 (N345, N319, N86);
nand NAND2_115 (N346, N319, N99);
nand NAND2_116 (N347, N319, N112);
nand NAND2_117 (N348, N330, N300);
nand NAND2_118 (N349, N331, N301);
nand NAND2_119 (N350, N332, N302);
nand NAND2_120 (N351, N333, N303);
nand NAND2_121 (N352, N335, N304);
nand NAND2_122 (N353, N337, N305);
nand NAND2_123 (N354, N339, N306);
nand NAND2_124 (N355, N341, N307);
nand NAND2_125 (N356, N343, N308);
  and AND9_126 (keyinput_Wire_0[22], N348, N349, N350, N351, N352, N353, N354, N355, N356);
  xnor keyGate_0_22(N357, keyinput22, keyinput_Wire_0[22]);
  not NOT1_127 (keyinput_Wire_0[23], N357);
  xnor keyGate_0_23(KeyNOTWire_0[13], keyinput23, keyinput_Wire_0[23]);
  not KeyNOTGate_0_13(N360, KeyNOTWire_0[13]);
not NOT1_128 (N370, N357);
nand NAND2_129 (N371, N14, N360);
nand NAND2_130 (N372, N360, N27);
nand NAND2_131 (N373, N360, N40);
nand NAND2_132 (N374, N360, N53);
nand NAND2_133 (N375, N360, N66);
nand NAND2_134 (N376, N360, N79);
nand NAND2_135 (N377, N360, N92);
nand NAND2_136 (N378, N360, N105);
nand NAND2_137 (N379, N360, N115);
nand NAND4_138 (N380, N4, N242, N334, N371);
nand NAND4_139 (N381, N246, N336, N372, N17);
nand NAND4_140 (N386, N250, N338, N373, N30);
  nand NAND4_141 (keyinput_Wire_0[24], N254, N340, N374, N43);
  xor keyGate_0_24(N393, keyinput24, keyinput_Wire_0[24]);
nand NAND4_142 (N399, N255, N342, N375, N56);
nand NAND4_143 (N404, N256, N344, N376, N69);
nand NAND4_144 (N407, N257, N345, N377, N82);
nand NAND4_145 (N411, N258, N346, N378, N95);
nand NAND4_146 (N414, N259, N347, N379, N108);
not NOT1_147 (N415, N380);
  and AND8_148 (keyinput_Wire_0[25], N381, N386, N393, N399, N404, N407, N411, N414);
  xnor keyGate_0_25(N416, keyinput25, keyinput_Wire_0[25]);
not NOT1_149 (N417, N393);
not NOT1_150 (N418, N404);
not NOT1_151 (N419, N407);
not NOT1_152 (N420, N411);
  nor NOR2_153 (keyinput_Wire_0[26], N415, N416);
  xnor keyGate_0_26(N421, keyinput26, keyinput_Wire_0[26]);
nand NAND2_154 (N422, N386, N417);
  nand NAND4_155 (keyinput_Wire_0[27], N386, N393, N418, N399);
  xor keyGate_0_27(KeyNOTWire_0[14], keyinput27, keyinput_Wire_0[27]);
  not KeyNOTGate_0_14(N425, KeyNOTWire_0[14]);
nand NAND3_156 (N428, N399, N393, N419);
  nand NAND4_157 (keyinput_Wire_0[28], N386, N393, N407, N420);
  xnor keyGate_0_28(KeyNOTWire_0[15], keyinput28, keyinput_Wire_0[28]);
  not KeyNOTGate_0_15(N429, KeyNOTWire_0[15]);
  nand NAND4_158 (keyinput_Wire_0[29], N381, N386, N422, N399);
  xnor keyGate_0_29(KeyNOTWire_0[16], keyinput29, keyinput_Wire_0[29]);
  not KeyNOTGate_0_16(N430, KeyNOTWire_0[16]);
  nand NAND4_159 (keyinput_Wire_0[30], N381, N386, N425, N428);
  xnor keyGate_0_30(KeyWire_0_1, keyinput30, keyinput_Wire_0[30]);
  xor flip_it (N431, KeyWire_0_1, KeyWire_0_2 );
  nand NAND4_160 (keyinput_Wire_0[31], N381, N422, N425, N429);
  xor keyGate_0_31(KeyNOTWire_0[17], keyinput31, keyinput_Wire_0[31]);
  not KeyNOTGate_0_17(N432, KeyNOTWire_0[17]);

AntiSAT some_name( KeyWire_0_2, N40, N89, N11, N56, N47, N21, N99, N43, N112, N8, N108, N50, N63, N95, N79, N69, N115, N60, N17, N37, N105, N14, N66, N86, N1, N102, N76, N4, N24, N27, N92, N53, N82, N34, N30, N73, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
       keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
       keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
       keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
       keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
       keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
       keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
       keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
       keyinput139);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N40, N89, N11, N56, N47, N21, N99, N43, N112, N8, N108, N50, N63, N95, N79, N69, N115, N60, N17, N37, N105, N14, N66, N86, N1, N102, N76, N4, N24, N27, N92, N53, N82, N34, N30, N73, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103 ,
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
        keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
        keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
        keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
        keyinput139);

  input keyinput104, keyinput105, keyinput106, keyinput107, keyinput108;
  input keyinput109, keyinput110, keyinput111, keyinput112, keyinput113;
  input keyinput114, keyinput115, keyinput116, keyinput117, keyinput118;
  input keyinput119, keyinput120, keyinput121, keyinput122, keyinput123;
  input keyinput124, keyinput125, keyinput126, keyinput127, keyinput128;
  input keyinput129, keyinput130, keyinput131, keyinput132, keyinput133;
  input keyinput134, keyinput135, keyinput136, keyinput137, keyinput138;
  input keyinput139;

  wire [0:35] keyNTin_Wire_1;
  wire [0:16] KeyNOTWire_1;

  input N40, N89, N11, N56, N47, N21, N99, N43, N112, N8, N108, N50, N63, N95, N79, N69, N115, N60, N17, N37, N105, N14, N66, N86, N1, N102, N76, N4, N24, N27, N92, N53, N82, N34, N30, N73;
  input keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73 ;

  xor  KeyGate0 (keyNTin_Wire_1[0], N40, keyinput32);
  xnor keyNTinGate_1_0(newWire_0, keyinput104, keyNTin_Wire_1[0]);
  xnor KeyGate1 (keyNTin_Wire_1[1], N89, keyinput33);
  xor keyNTinGate_1_1(newWire_1, keyinput105, keyNTin_Wire_1[1]);
  xnor KeyGate2 (newWire_2, N11, keyinput34);
  xor  KeyGate3 (keyNTin_Wire_1[2], N56, keyinput35);
  xnor keyNTinGate_1_2(KeyNOTWire_1[0], keyinput106, keyNTin_Wire_1[2]);
  not KeyNOTGate_1_0(newWire_3, KeyNOTWire_1[0]);
  xnor KeyGate4 (keyNTin_Wire_1[3], N47, keyinput36);
  xnor keyNTinGate_1_3(newWire_4, keyinput107, keyNTin_Wire_1[3]);
  xnor KeyGate5 (newWire_5, N21, keyinput37);
  xor  KeyGate6 (newWire_6, N99, keyinput38);
  xor  KeyGate7 (keyNTin_Wire_1[4], N43, keyinput39);
  xnor keyNTinGate_1_4(newWire_7, keyinput108, keyNTin_Wire_1[4]);
  xor  KeyGate8 (newWire_8, N112, keyinput40);
  xnor KeyGate9 (newWire_9, N8, keyinput41);
  xor  KeyGate10 (keyNTin_Wire_1[5], N108, keyinput42);
  xnor keyNTinGate_1_5(newWire_10, keyinput109, keyNTin_Wire_1[5]);
  xnor KeyGate11 (keyNTin_Wire_1[6], N50, keyinput43);
  xor keyNTinGate_1_6(KeyNOTWire_1[1], keyinput110, keyNTin_Wire_1[6]);
  not KeyNOTGate_1_1(newWire_11, KeyNOTWire_1[1]);
  xor  KeyGate12 (keyNTin_Wire_1[7], N63, keyinput44);
  xor keyNTinGate_1_7(KeyNOTWire_1[2], keyinput111, keyNTin_Wire_1[7]);
  not KeyNOTGate_1_2(newWire_12, KeyNOTWire_1[2]);
  xor  KeyGate13 (newWire_13, N95, keyinput45);
  xor  KeyGate14 (newWire_14, N79, keyinput46);
  xnor KeyGate15 (newWire_15, N69, keyinput47);
  xnor KeyGate16 (keyNTin_Wire_1[8], N115, keyinput48);
  xor keyNTinGate_1_8(newWire_16, keyinput112, keyNTin_Wire_1[8]);
  xnor KeyGate17 (newWire_17, N60, keyinput49);
  xnor KeyGate18 (keyNTin_Wire_1[9], N17, keyinput50);
  xor keyNTinGate_1_9(KeyNOTWire_1[3], keyinput113, keyNTin_Wire_1[9]);
  not KeyNOTGate_1_3(newWire_18, KeyNOTWire_1[3]);
  xor  KeyGate19 (keyNTin_Wire_1[10], N37, keyinput51);
  xor keyNTinGate_1_10(newWire_19, keyinput114, keyNTin_Wire_1[10]);
  xnor KeyGate20 (newWire_20, N105, keyinput52);
  xnor KeyGate21 (keyNTin_Wire_1[11], N14, keyinput53);
  xor keyNTinGate_1_11(KeyNOTWire_1[4], keyinput115, keyNTin_Wire_1[11]);
  not KeyNOTGate_1_4(newWire_21, KeyNOTWire_1[4]);
  xnor KeyGate22 (keyNTin_Wire_1[12], N66, keyinput54);
  xor keyNTinGate_1_12(KeyNOTWire_1[5], keyinput116, keyNTin_Wire_1[12]);
  not KeyNOTGate_1_5(newWire_22, KeyNOTWire_1[5]);
  xor  KeyGate23 (keyNTin_Wire_1[13], N86, keyinput55);
  xor keyNTinGate_1_13(KeyNOTWire_1[6], keyinput117, keyNTin_Wire_1[13]);
  not KeyNOTGate_1_6(newWire_23, KeyNOTWire_1[6]);
  xnor KeyGate24 (keyNTin_Wire_1[14], N1, keyinput56);
  xor keyNTinGate_1_14(KeyNOTWire_1[7], keyinput118, keyNTin_Wire_1[14]);
  not KeyNOTGate_1_7(newWire_24, KeyNOTWire_1[7]);
  xnor KeyGate25 (keyNTin_Wire_1[15], N102, keyinput57);
  xnor keyNTinGate_1_15(newWire_25, keyinput119, keyNTin_Wire_1[15]);
  xnor KeyGate26 (newWire_26, N76, keyinput58);
  xor  KeyGate27 (newWire_27, N4, keyinput59);
  xor  KeyGate28 (keyNTin_Wire_1[16], N24, keyinput60);
  xnor keyNTinGate_1_16(KeyNOTWire_1[8], keyinput120, keyNTin_Wire_1[16]);
  not KeyNOTGate_1_8(newWire_28, KeyNOTWire_1[8]);
  xor  KeyGate29 (keyNTin_Wire_1[17], N27, keyinput61);
  xnor keyNTinGate_1_17(newWire_29, keyinput121, keyNTin_Wire_1[17]);
  xor  KeyGate30 (newWire_30, N92, keyinput62);
  xor  KeyGate31 (newWire_31, N53, keyinput63);
  xnor KeyGate32 (newWire_32, N82, keyinput64);
  xor  KeyGate33 (keyNTin_Wire_1[18], N34, keyinput65);
  xor keyNTinGate_1_18(KeyNOTWire_1[9], keyinput122, keyNTin_Wire_1[18]);
  not KeyNOTGate_1_9(newWire_33, KeyNOTWire_1[9]);
  xor  KeyGate34 (keyNTin_Wire_1[19], N30, keyinput66);
  xnor keyNTinGate_1_19(newWire_34, keyinput123, keyNTin_Wire_1[19]);
  xnor KeyGate35 (keyNTin_Wire_1[20], N73, keyinput67);
  xor keyNTinGate_1_20(newWire_35, keyinput124, keyNTin_Wire_1[20]);
  xnor KeyGate36 (newWire_36, N40, keyinput68);
  xor  KeyGate37 (keyNTin_Wire_1[21], N89, keyinput69);
  xnor keyNTinGate_1_21(newWire_37, keyinput125, keyNTin_Wire_1[21]);
  xor  KeyGate38 (newWire_38, N11, keyinput70);
  xor  KeyGate39 (newWire_39, N56, keyinput71);
  xnor KeyGate40 (keyNTin_Wire_1[22], N47, keyinput72);
  xor keyNTinGate_1_22(newWire_40, keyinput126, keyNTin_Wire_1[22]);
  xnor KeyGate41 (newWire_41, N21, keyinput73);
  xor  KeyGate42 (keyNTin_Wire_1[23], N99, keyinput74);
  xnor keyNTinGate_1_23(KeyNOTWire_1[10], keyinput127, keyNTin_Wire_1[23]);
  not KeyNOTGate_1_10(newWire_42, KeyNOTWire_1[10]);
  xnor KeyGate43 (newWire_43, N43, keyinput75);
  xor  KeyGate44 (newWire_44, N112, keyinput76);
  xor  KeyGate45 (newWire_45, N8, keyinput77);
  xnor KeyGate46 (newWire_46, N108, keyinput78);
  xnor KeyGate47 (keyNTin_Wire_1[24], N50, keyinput79);
  xor keyNTinGate_1_24(newWire_47, keyinput128, keyNTin_Wire_1[24]);
  xor  KeyGate48 (newWire_48, N63, keyinput80);
  xnor KeyGate49 (newWire_49, N95, keyinput81);
  xnor KeyGate50 (newWire_50, N79, keyinput82);
  xor  KeyGate51 (keyNTin_Wire_1[25], N69, keyinput83);
  xnor keyNTinGate_1_25(KeyNOTWire_1[11], keyinput129, keyNTin_Wire_1[25]);
  not KeyNOTGate_1_11(newWire_51, KeyNOTWire_1[11]);
  xnor KeyGate52 (keyNTin_Wire_1[26], N115, keyinput84);
  xor keyNTinGate_1_26(newWire_52, keyinput130, keyNTin_Wire_1[26]);
  xnor KeyGate53 (newWire_53, N60, keyinput85);
  xnor KeyGate54 (newWire_54, N17, keyinput86);
  xor  KeyGate55 (newWire_55, N37, keyinput87);
  xnor KeyGate56 (newWire_56, N105, keyinput88);
  xor  KeyGate57 (newWire_57, N14, keyinput89);
  xnor KeyGate58 (keyNTin_Wire_1[27], N66, keyinput90);
  xnor keyNTinGate_1_27(newWire_58, keyinput131, keyNTin_Wire_1[27]);
  xnor KeyGate59 (newWire_59, N86, keyinput91);
  xor  KeyGate60 (newWire_60, N1, keyinput92);
  xnor KeyGate61 (newWire_61, N102, keyinput93);
  xnor KeyGate62 (keyNTin_Wire_1[28], N76, keyinput94);
  xnor keyNTinGate_1_28(KeyNOTWire_1[12], keyinput132, keyNTin_Wire_1[28]);
  not KeyNOTGate_1_12(newWire_62, KeyNOTWire_1[12]);
  xnor KeyGate63 (keyNTin_Wire_1[29], N4, keyinput95);
  xnor keyNTinGate_1_29(KeyNOTWire_1[13], keyinput133, keyNTin_Wire_1[29]);
  not KeyNOTGate_1_13(newWire_63, KeyNOTWire_1[13]);
  xnor KeyGate64 (keyNTin_Wire_1[30], N24, keyinput96);
  xor keyNTinGate_1_30(KeyNOTWire_1[14], keyinput134, keyNTin_Wire_1[30]);
  not KeyNOTGate_1_14(newWire_64, KeyNOTWire_1[14]);
  xor  KeyGate65 (keyNTin_Wire_1[31], N27, keyinput97);
  xor keyNTinGate_1_31(newWire_65, keyinput135, keyNTin_Wire_1[31]);
  xnor KeyGate66 (newWire_66, N92, keyinput98);
  xnor KeyGate67 (newWire_67, N53, keyinput99);
  xor  KeyGate68 (newWire_68, N82, keyinput100);
  xnor KeyGate69 (newWire_69, N34, keyinput101);
  xor  KeyGate70 (keyNTin_Wire_1[32], N30, keyinput102);
  xnor keyNTinGate_1_32(KeyNOTWire_1[15], keyinput136, keyNTin_Wire_1[32]);
  not KeyNOTGate_1_15(newWire_70, KeyNOTWire_1[15]);
  xnor KeyGate71 (keyNTin_Wire_1[33], N73, keyinput103);
  xor keyNTinGate_1_33(KeyNOTWire_1[16], keyinput137, keyNTin_Wire_1[33]);
  not KeyNOTGate_1_16(newWire_71, KeyNOTWire_1[16]);
  and some_function (keyNTin_Wire_1[34], newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35 );
  xor keyNTinGate_1_34(newWire_72, keyinput138, keyNTin_Wire_1[34]);
  nand compl_function (newWire_73, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71);
  and finalAND (keyNTin_Wire_1[35], newWire_72, newWire_73);
  xor keyNTinGate_1_35(KeyWire_0_2, keyinput139, keyNTin_Wire_1[35]);

endmodule /* AntiSAT */
