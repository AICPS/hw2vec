`timescale 1ns / 1ps
module top (G1,G10,G11,G12,G13,G1324,G1325,G1326,G1327,G1328,G1329,G1330,
  G1331,G1332,G1333,G1334,G1335,G1336,G1337,G1338,G1339,G1340,G1341,G1342,
  G1343,G1344,G1345,G1346,G1347,G1348,G1349,G1350,G1351,G1352,G1353,G1354,
  G1355,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G3,
                  G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G4,G40,G41,G5,G6,G7,G8,G9,
        keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4,
        keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9,
        keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14,
        keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19,
        keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24,
        keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29,
        keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34,
        keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39,
        keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44,
        keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49,
        keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54,
        keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59,
        keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64,
        keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69,
        keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74,
        keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79,
        keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84,
        keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89,
        keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94,
        keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99,
        keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104,
        keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109,
        keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114,
        keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119,
        keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124,
        keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129,
        keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134,
        keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139,
        keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144,
        keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149,
        keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154,
        keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159,
        keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164,
        keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169,
        keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174,
        keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179,
        keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184,
        keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189,
        keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194,
        keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199,
        keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204,
        keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209,
        keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214,
        keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219,
        keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224,
        keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229,
        keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234,
        keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239,
        keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244,
        keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249,
        keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254,
        keyIn_0_255);

  input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4;
  input keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9;
  input keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14;
  input keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19;
  input keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24;
  input keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29;
  input keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34;
  input keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39;
  input keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44;
  input keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49;
  input keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54;
  input keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59;
  input keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64;
  input keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69;
  input keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74;
  input keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79;
  input keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84;
  input keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89;
  input keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94;
  input keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99;
  input keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104;
  input keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109;
  input keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114;
  input keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119;
  input keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124;
  input keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129;
  input keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134;
  input keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139;
  input keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144;
  input keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149;
  input keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154;
  input keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159;
  input keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164;
  input keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169;
  input keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174;
  input keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179;
  input keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184;
  input keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189;
  input keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194;
  input keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199;
  input keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204;
  input keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209;
  input keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214;
  input keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219;
  input keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224;
  input keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229;
  input keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234;
  input keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239;
  input keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244;
  input keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249;
  input keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254;
  input keyIn_0_255;

  wire [0:255] KeyWire_0;
  wire [0:137] KeyNOTWire_0;
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
  G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,
  G40,G41;
output G1324,G1325,G1326,G1327,G1328,G1329,G1330,G1331,G1332,G1333,G1334,G1335,
  G1336,G1337,G1338,G1339,G1340,G1341,G1342,G1343,G1344,G1345,G1346,G1347,
  G1348,G1349,G1350,G1351,G1352,G1353,G1354,G1355;

  wire G242,G245,G248,G251,G254,G257,G260,G263,G266,G269,G272,G275,G278,G281,
    G284,G287,G290,G293,G296,G299,G302,G305,G308,G311,G314,G317,G320,G323,G326,
    G329,G332,G335,G338,G341,G344,G347,G350,G353,G356,G359,G362,G363,G364,G365,
    G366,G367,G368,G369,G370,G371,G372,G373,G374,G375,G376,G377,G378,G379,G380,
    G381,G382,G383,G384,G385,G386,G387,G388,G389,G390,G391,G392,G393,G394,G395,
    G396,G397,G398,G399,G400,G401,G402,G403,G404,G405,G406,G407,G408,G409,G410,
    G411,G412,G413,G414,G415,G416,G417,G418,G419,G420,G421,G422,G423,G424,G425,
    G426,G429,G432,G435,G438,G441,G444,G447,G450,G453,G456,G459,G462,G465,G468,
    G471,G474,G477,G480,G483,G486,G489,G492,G495,G498,G501,G504,G507,G510,G513,
    G516,G519,G522,G525,G528,G531,G534,G537,G540,G543,G546,G549,G552,G555,G558,
    G561,G564,G567,G570,G571,G572,G573,G574,G575,G576,G577,G578,G579,G580,G581,
    G582,G583,G584,G585,G586,G587,G588,G589,G590,G591,G592,G593,G594,G595,G596,
    G597,G598,G599,G600,G601,G602,G607,G612,G617,G622,G627,G632,G637,G642,G645,
    G648,G651,G654,G657,G660,G663,G666,G669,G672,G675,G678,G681,G684,G687,G690,
    G691,G692,G693,G694,G695,G696,G697,G698,G699,G700,G701,G702,G703,G704,G705,
    G706,G709,G712,G715,G718,G721,G724,G727,G730,G733,G736,G739,G742,G745,G748,
    G751,G754,G755,G756,G757,G758,G759,G760,G761,G762,G763,G764,G765,G766,G767,
    G768,G769,G770,G773,G776,G779,G782,G785,G788,G791,G794,G797,G800,G803,G806,
    G809,G812,G815,G818,G819,G820,G821,G822,G823,G824,G825,G826,G827,G828,G829,
    G830,G831,G832,G833,G834,G847,G860,G873,G886,G899,G912,G925,G938,G939,G940,
    G941,G942,G943,G944,G945,G946,G947,G948,G949,G950,G951,G952,G953,G954,G955,
    G956,G957,G958,G959,G960,G961,G962,G963,G964,G965,G966,G967,G968,G969,G970,
    G971,G972,G973,G974,G975,G976,G977,G978,G979,G980,G981,G982,G983,G984,G985,
    G986,G991,G996,G1001,G1006,G1011,G1016,G1021,G1026,G1031,G1036,G1039,G1042,
    G1045,G1048,G1051,G1054,G1057,G1060,G1063,G1066,G1069,G1072,G1075,G1078,
    G1081,G1084,G1087,G1090,G1093,G1096,G1099,G1102,G1105,G1108,G1111,G1114,
    G1117,G1120,G1123,G1126,G1129,G1132,G1135,G1138,G1141,G1144,G1147,G1150,
    G1153,G1156,G1159,G1162,G1165,G1168,G1171,G1174,G1177,G1180,G1183,G1186,
    G1189,G1192,G1195,G1198,G1201,G1204,G1207,G1210,G1213,G1216,G1219,G1222,
    G1225,G1228,G1229,G1230,G1231,G1232,G1233,G1234,G1235,G1236,G1237,G1238,
    G1239,G1240,G1241,G1242,G1243,G1244,G1245,G1246,G1247,G1248,G1249,G1250,
    G1251,G1252,G1253,G1254,G1255,G1256,G1257,G1258,G1259,G1260,G1261,G1262,
    G1263,G1264,G1265,G1266,G1267,G1268,G1269,G1270,G1271,G1272,G1273,G1274,
    G1275,G1276,G1277,G1278,G1279,G1280,G1281,G1282,G1283,G1284,G1285,G1286,
    G1287,G1288,G1289,G1290,G1291,G1292,G1293,G1294,G1295,G1296,G1297,G1298,
    G1299,G1300,G1301,G1302,G1303,G1304,G1305,G1306,G1307,G1308,G1309,G1310,
    G1311,G1312,G1313,G1314,G1315,G1316,G1317,G1318,G1319,G1320,G1321,G1322,
    G1323;

  and AND2_0(G242,G33,G41);
  and AND2_1(G245,G34,G41);
  and AND2_2(KeyWire_0[0], G35,G41);
  xnor KeyGate_0_0(KeyNOTWire_0[0], keyIn_0_0, KeyWire_0[0]);
  not KeyNOTGate_0_0(G248, KeyNOTWire_0[0]);
  and AND2_3(KeyWire_0[1], G36,G41);
  xnor KeyGate_0_1(KeyNOTWire_0[1], keyIn_0_1, KeyWire_0[1]);
  not KeyNOTGate_0_1(G251, KeyNOTWire_0[1]);
  and AND2_4(G254,G37,G41);
  and AND2_5(G257,G38,G41);
  and AND2_6(KeyWire_0[2], G39,G41);
  xnor KeyGate_0_2(G260, keyIn_0_2, KeyWire_0[2]);
  and AND2_7(G263,G40,G41);
  nand NAND2_0(KeyWire_0[3], G1,G2);
  xnor KeyGate_0_3(KeyNOTWire_0[2], keyIn_0_3, KeyWire_0[3]);
  not KeyNOTGate_0_2(G266, KeyNOTWire_0[2]);
  nand NAND2_1(G269,G3,G4);
  nand NAND2_2(G272,G5,G6);
  nand NAND2_3(G275,G7,G8);
  nand NAND2_4(KeyWire_0[4], G9,G10);
  xor KeyGate_0_4(G278, keyIn_0_4, KeyWire_0[4]);
  nand NAND2_5(G281,G11,G12);
  nand NAND2_6(KeyWire_0[5], G13,G14);
  xnor KeyGate_0_5(G284, keyIn_0_5, KeyWire_0[5]);
  nand NAND2_7(G287,G15,G16);
  nand NAND2_8(KeyWire_0[6], G17,G18);
  xnor KeyGate_0_6(KeyNOTWire_0[3], keyIn_0_6, KeyWire_0[6]);
  not KeyNOTGate_0_3(G290, KeyNOTWire_0[3]);
  nand NAND2_9(KeyWire_0[7], G19,G20);
  xnor KeyGate_0_7(KeyNOTWire_0[4], keyIn_0_7, KeyWire_0[7]);
  not KeyNOTGate_0_4(G293, KeyNOTWire_0[4]);
  nand NAND2_10(KeyWire_0[8], G21,G22);
  xor KeyGate_0_8(KeyNOTWire_0[5], keyIn_0_8, KeyWire_0[8]);
  not KeyNOTGate_0_5(G296, KeyNOTWire_0[5]);
  nand NAND2_11(G299,G23,G24);
  nand NAND2_12(KeyWire_0[9], G25,G26);
  xor KeyGate_0_9(G302, keyIn_0_9, KeyWire_0[9]);
  nand NAND2_13(G305,G27,G28);
  nand NAND2_14(KeyWire_0[10], G29,G30);
  xor KeyGate_0_10(G308, keyIn_0_10, KeyWire_0[10]);
  nand NAND2_15(KeyWire_0[11], G31,G32);
  xnor KeyGate_0_11(KeyNOTWire_0[6], keyIn_0_11, KeyWire_0[11]);
  not KeyNOTGate_0_6(G311, KeyNOTWire_0[6]);
  nand NAND2_16(G314,G1,G5);
  nand NAND2_17(KeyWire_0[12], G9,G13);
  xor KeyGate_0_12(G317, keyIn_0_12, KeyWire_0[12]);
  nand NAND2_18(G320,G2,G6);
  nand NAND2_19(G323,G10,G14);
  nand NAND2_20(G326,G3,G7);
  nand NAND2_21(G329,G11,G15);
  nand NAND2_22(G332,G4,G8);
  nand NAND2_23(G335,G12,G16);
  nand NAND2_24(KeyWire_0[13], G17,G21);
  xor KeyGate_0_13(KeyNOTWire_0[7], keyIn_0_13, KeyWire_0[13]);
  not KeyNOTGate_0_7(G338, KeyNOTWire_0[7]);
  nand NAND2_25(KeyWire_0[14], G25,G29);
  xnor KeyGate_0_14(G341, keyIn_0_14, KeyWire_0[14]);
  nand NAND2_26(KeyWire_0[15], G18,G22);
  xor KeyGate_0_15(G344, keyIn_0_15, KeyWire_0[15]);
  nand NAND2_27(G347,G26,G30);
  nand NAND2_28(KeyWire_0[16], G19,G23);
  xnor KeyGate_0_16(KeyNOTWire_0[8], keyIn_0_16, KeyWire_0[16]);
  not KeyNOTGate_0_8(G350, KeyNOTWire_0[8]);
  nand NAND2_29(KeyWire_0[17], G27,G31);
  xor KeyGate_0_17(G353, keyIn_0_17, KeyWire_0[17]);
  nand NAND2_30(G356,G20,G24);
  nand NAND2_31(KeyWire_0[18], G28,G32);
  xor KeyGate_0_18(KeyNOTWire_0[9], keyIn_0_18, KeyWire_0[18]);
  not KeyNOTGate_0_9(G359, KeyNOTWire_0[9]);
  nand NAND2_32(G362,G1,G266);
  nand NAND2_33(KeyWire_0[19], G2,G266);
  xor KeyGate_0_19(KeyNOTWire_0[10], keyIn_0_19, KeyWire_0[19]);
  not KeyNOTGate_0_10(G363, KeyNOTWire_0[10]);
  nand NAND2_34(KeyWire_0[20], G3,G269);
  xor KeyGate_0_20(KeyNOTWire_0[11], keyIn_0_20, KeyWire_0[20]);
  not KeyNOTGate_0_11(G364, KeyNOTWire_0[11]);
  nand NAND2_35(G365,G4,G269);
  nand NAND2_36(G366,G5,G272);
  nand NAND2_37(G367,G6,G272);
  nand NAND2_38(G368,G7,G275);
  nand NAND2_39(KeyWire_0[21], G8,G275);
  xnor KeyGate_0_21(KeyNOTWire_0[12], keyIn_0_21, KeyWire_0[21]);
  not KeyNOTGate_0_12(G369, KeyNOTWire_0[12]);
  nand NAND2_40(G370,G9,G278);
  nand NAND2_41(KeyWire_0[22], G10,G278);
  xnor KeyGate_0_22(G371, keyIn_0_22, KeyWire_0[22]);
  nand NAND2_42(G372,G11,G281);
  nand NAND2_43(G373,G12,G281);
  nand NAND2_44(KeyWire_0[23], G13,G284);
  xnor KeyGate_0_23(G374, keyIn_0_23, KeyWire_0[23]);
  nand NAND2_45(KeyWire_0[24], G14,G284);
  xnor KeyGate_0_24(KeyNOTWire_0[13], keyIn_0_24, KeyWire_0[24]);
  not KeyNOTGate_0_13(G375, KeyNOTWire_0[13]);
  nand NAND2_46(KeyWire_0[25], G15,G287);
  xnor KeyGate_0_25(G376, keyIn_0_25, KeyWire_0[25]);
  nand NAND2_47(KeyWire_0[26], G16,G287);
  xor KeyGate_0_26(G377, keyIn_0_26, KeyWire_0[26]);
  nand NAND2_48(G378,G17,G290);
  nand NAND2_49(G379,G18,G290);
  nand NAND2_50(G380,G19,G293);
  nand NAND2_51(KeyWire_0[27], G20,G293);
  xnor KeyGate_0_27(G381, keyIn_0_27, KeyWire_0[27]);
  nand NAND2_52(G382,G21,G296);
  nand NAND2_53(KeyWire_0[28], G22,G296);
  xor KeyGate_0_28(KeyNOTWire_0[14], keyIn_0_28, KeyWire_0[28]);
  not KeyNOTGate_0_14(G383, KeyNOTWire_0[14]);
  nand NAND2_54(G384,G23,G299);
  nand NAND2_55(G385,G24,G299);
  nand NAND2_56(G386,G25,G302);
  nand NAND2_57(G387,G26,G302);
  nand NAND2_58(G388,G27,G305);
  nand NAND2_59(KeyWire_0[29], G28,G305);
  xnor KeyGate_0_29(KeyNOTWire_0[15], keyIn_0_29, KeyWire_0[29]);
  not KeyNOTGate_0_15(G389, KeyNOTWire_0[15]);
  nand NAND2_60(G390,G29,G308);
  nand NAND2_61(G391,G30,G308);
  nand NAND2_62(G392,G31,G311);
  nand NAND2_63(G393,G32,G311);
  nand NAND2_64(KeyWire_0[30], G1,G314);
  xnor KeyGate_0_30(G394, keyIn_0_30, KeyWire_0[30]);
  nand NAND2_65(KeyWire_0[31], G5,G314);
  xnor KeyGate_0_31(KeyNOTWire_0[16], keyIn_0_31, KeyWire_0[31]);
  not KeyNOTGate_0_16(G395, KeyNOTWire_0[16]);
  nand NAND2_66(G396,G9,G317);
  nand NAND2_67(G397,G13,G317);
  nand NAND2_68(G398,G2,G320);
  nand NAND2_69(G399,G6,G320);
  nand NAND2_70(G400,G10,G323);
  nand NAND2_71(KeyWire_0[32], G14,G323);
  xor KeyGate_0_32(G401, keyIn_0_32, KeyWire_0[32]);
  nand NAND2_72(G402,G3,G326);
  nand NAND2_73(KeyWire_0[33], G7,G326);
  xor KeyGate_0_33(G403, keyIn_0_33, KeyWire_0[33]);
  nand NAND2_74(G404,G11,G329);
  nand NAND2_75(G405,G15,G329);
  nand NAND2_76(KeyWire_0[34], G4,G332);
  xor KeyGate_0_34(G406, keyIn_0_34, KeyWire_0[34]);
  nand NAND2_77(G407,G8,G332);
  nand NAND2_78(KeyWire_0[35], G12,G335);
  xnor KeyGate_0_35(G408, keyIn_0_35, KeyWire_0[35]);
  nand NAND2_79(KeyWire_0[36], G16,G335);
  xor KeyGate_0_36(G409, keyIn_0_36, KeyWire_0[36]);
  nand NAND2_80(KeyWire_0[37], G17,G338);
  xnor KeyGate_0_37(KeyNOTWire_0[17], keyIn_0_37, KeyWire_0[37]);
  not KeyNOTGate_0_17(G410, KeyNOTWire_0[17]);
  nand NAND2_81(KeyWire_0[38], G21,G338);
  xnor KeyGate_0_38(KeyNOTWire_0[18], keyIn_0_38, KeyWire_0[38]);
  not KeyNOTGate_0_18(G411, KeyNOTWire_0[18]);
  nand NAND2_82(KeyWire_0[39], G25,G341);
  xor KeyGate_0_39(KeyNOTWire_0[19], keyIn_0_39, KeyWire_0[39]);
  not KeyNOTGate_0_19(G412, KeyNOTWire_0[19]);
  nand NAND2_83(G413,G29,G341);
  nand NAND2_84(KeyWire_0[40], G18,G344);
  xor KeyGate_0_40(G414, keyIn_0_40, KeyWire_0[40]);
  nand NAND2_85(G415,G22,G344);
  nand NAND2_86(G416,G26,G347);
  nand NAND2_87(KeyWire_0[41], G30,G347);
  xnor KeyGate_0_41(KeyNOTWire_0[20], keyIn_0_41, KeyWire_0[41]);
  not KeyNOTGate_0_20(G417, KeyNOTWire_0[20]);
  nand NAND2_88(G418,G19,G350);
  nand NAND2_89(G419,G23,G350);
  nand NAND2_90(KeyWire_0[42], G27,G353);
  xnor KeyGate_0_42(KeyNOTWire_0[21], keyIn_0_42, KeyWire_0[42]);
  not KeyNOTGate_0_21(G420, KeyNOTWire_0[21]);
  nand NAND2_91(G421,G31,G353);
  nand NAND2_92(KeyWire_0[43], G20,G356);
  xor KeyGate_0_43(KeyNOTWire_0[22], keyIn_0_43, KeyWire_0[43]);
  not KeyNOTGate_0_22(G422, KeyNOTWire_0[22]);
  nand NAND2_93(G423,G24,G356);
  nand NAND2_94(KeyWire_0[44], G28,G359);
  xor KeyGate_0_44(KeyNOTWire_0[23], keyIn_0_44, KeyWire_0[44]);
  not KeyNOTGate_0_23(G424, KeyNOTWire_0[23]);
  nand NAND2_95(KeyWire_0[45], G32,G359);
  xor KeyGate_0_45(KeyNOTWire_0[24], keyIn_0_45, KeyWire_0[45]);
  not KeyNOTGate_0_24(G425, KeyNOTWire_0[24]);
  nand NAND2_96(G426,G362,G363);
  nand NAND2_97(KeyWire_0[46], G364,G365);
  xor KeyGate_0_46(KeyNOTWire_0[25], keyIn_0_46, KeyWire_0[46]);
  not KeyNOTGate_0_25(G429, KeyNOTWire_0[25]);
  nand NAND2_98(G432,G366,G367);
  nand NAND2_99(KeyWire_0[47], G368,G369);
  xor KeyGate_0_47(G435, keyIn_0_47, KeyWire_0[47]);
  nand NAND2_100(KeyWire_0[48], G370,G371);
  xor KeyGate_0_48(G438, keyIn_0_48, KeyWire_0[48]);
  nand NAND2_101(KeyWire_0[49], G372,G373);
  xor KeyGate_0_49(KeyNOTWire_0[26], keyIn_0_49, KeyWire_0[49]);
  not KeyNOTGate_0_26(G441, KeyNOTWire_0[26]);
  nand NAND2_102(KeyWire_0[50], G374,G375);
  xor KeyGate_0_50(G444, keyIn_0_50, KeyWire_0[50]);
  nand NAND2_103(KeyWire_0[51], G376,G377);
  xor KeyGate_0_51(G447, keyIn_0_51, KeyWire_0[51]);
  nand NAND2_104(KeyWire_0[52], G378,G379);
  xor KeyGate_0_52(KeyNOTWire_0[27], keyIn_0_52, KeyWire_0[52]);
  not KeyNOTGate_0_27(G450, KeyNOTWire_0[27]);
  nand NAND2_105(KeyWire_0[53], G380,G381);
  xnor KeyGate_0_53(KeyNOTWire_0[28], keyIn_0_53, KeyWire_0[53]);
  not KeyNOTGate_0_28(G453, KeyNOTWire_0[28]);
  nand NAND2_106(KeyWire_0[54], G382,G383);
  xor KeyGate_0_54(KeyNOTWire_0[29], keyIn_0_54, KeyWire_0[54]);
  not KeyNOTGate_0_29(G456, KeyNOTWire_0[29]);
  nand NAND2_107(G459,G384,G385);
  nand NAND2_108(G462,G386,G387);
  nand NAND2_109(G465,G388,G389);
  nand NAND2_110(G468,G390,G391);
  nand NAND2_111(KeyWire_0[55], G392,G393);
  xor KeyGate_0_55(G471, keyIn_0_55, KeyWire_0[55]);
  nand NAND2_112(KeyWire_0[56], G394,G395);
  xnor KeyGate_0_56(G474, keyIn_0_56, KeyWire_0[56]);
  nand NAND2_113(KeyWire_0[57], G396,G397);
  xor KeyGate_0_57(KeyNOTWire_0[30], keyIn_0_57, KeyWire_0[57]);
  not KeyNOTGate_0_30(G477, KeyNOTWire_0[30]);
  nand NAND2_114(G480,G398,G399);
  nand NAND2_115(KeyWire_0[58], G400,G401);
  xor KeyGate_0_58(KeyNOTWire_0[31], keyIn_0_58, KeyWire_0[58]);
  not KeyNOTGate_0_31(G483, KeyNOTWire_0[31]);
  nand NAND2_116(G486,G402,G403);
  nand NAND2_117(G489,G404,G405);
  nand NAND2_118(KeyWire_0[59], G406,G407);
  xnor KeyGate_0_59(G492, keyIn_0_59, KeyWire_0[59]);
  nand NAND2_119(KeyWire_0[60], G408,G409);
  xnor KeyGate_0_60(KeyNOTWire_0[32], keyIn_0_60, KeyWire_0[60]);
  not KeyNOTGate_0_32(G495, KeyNOTWire_0[32]);
  nand NAND2_120(G498,G410,G411);
  nand NAND2_121(KeyWire_0[61], G412,G413);
  xnor KeyGate_0_61(KeyNOTWire_0[33], keyIn_0_61, KeyWire_0[61]);
  not KeyNOTGate_0_33(G501, KeyNOTWire_0[33]);
  nand NAND2_122(G504,G414,G415);
  nand NAND2_123(KeyWire_0[62], G416,G417);
  xnor KeyGate_0_62(KeyNOTWire_0[34], keyIn_0_62, KeyWire_0[62]);
  not KeyNOTGate_0_34(G507, KeyNOTWire_0[34]);
  nand NAND2_124(G510,G418,G419);
  nand NAND2_125(G513,G420,G421);
  nand NAND2_126(KeyWire_0[63], G422,G423);
  xnor KeyGate_0_63(G516, keyIn_0_63, KeyWire_0[63]);
  nand NAND2_127(G519,G424,G425);
  nand NAND2_128(G522,G426,G429);
  nand NAND2_129(G525,G432,G435);
  nand NAND2_130(G528,G438,G441);
  nand NAND2_131(KeyWire_0[64], G444,G447);
  xnor KeyGate_0_64(G531, keyIn_0_64, KeyWire_0[64]);
  nand NAND2_132(KeyWire_0[65], G450,G453);
  xnor KeyGate_0_65(G534, keyIn_0_65, KeyWire_0[65]);
  nand NAND2_133(G537,G456,G459);
  nand NAND2_134(G540,G462,G465);
  nand NAND2_135(G543,G468,G471);
  nand NAND2_136(KeyWire_0[66], G474,G477);
  xor KeyGate_0_66(G546, keyIn_0_66, KeyWire_0[66]);
  nand NAND2_137(KeyWire_0[67], G480,G483);
  xnor KeyGate_0_67(G549, keyIn_0_67, KeyWire_0[67]);
  nand NAND2_138(KeyWire_0[68], G486,G489);
  xnor KeyGate_0_68(KeyNOTWire_0[35], keyIn_0_68, KeyWire_0[68]);
  not KeyNOTGate_0_35(G552, KeyNOTWire_0[35]);
  nand NAND2_139(G555,G492,G495);
  nand NAND2_140(G558,G498,G501);
  nand NAND2_141(G561,G504,G507);
  nand NAND2_142(KeyWire_0[69], G510,G513);
  xnor KeyGate_0_69(KeyNOTWire_0[36], keyIn_0_69, KeyWire_0[69]);
  not KeyNOTGate_0_36(G564, KeyNOTWire_0[36]);
  nand NAND2_143(G567,G516,G519);
  nand NAND2_144(KeyWire_0[70], G426,G522);
  xor KeyGate_0_70(KeyNOTWire_0[37], keyIn_0_70, KeyWire_0[70]);
  not KeyNOTGate_0_37(G570, KeyNOTWire_0[37]);
  nand NAND2_145(G571,G429,G522);
  nand NAND2_146(G572,G432,G525);
  nand NAND2_147(G573,G435,G525);
  nand NAND2_148(KeyWire_0[71], G438,G528);
  xor KeyGate_0_71(G574, keyIn_0_71, KeyWire_0[71]);
  nand NAND2_149(G575,G441,G528);
  nand NAND2_150(KeyWire_0[72], G444,G531);
  xnor KeyGate_0_72(G576, keyIn_0_72, KeyWire_0[72]);
  nand NAND2_151(KeyWire_0[73], G447,G531);
  xnor KeyGate_0_73(G577, keyIn_0_73, KeyWire_0[73]);
  nand NAND2_152(G578,G450,G534);
  nand NAND2_153(G579,G453,G534);
  nand NAND2_154(KeyWire_0[74], G456,G537);
  xnor KeyGate_0_74(KeyNOTWire_0[38], keyIn_0_74, KeyWire_0[74]);
  not KeyNOTGate_0_38(G580, KeyNOTWire_0[38]);
  nand NAND2_155(KeyWire_0[75], G459,G537);
  xor KeyGate_0_75(KeyNOTWire_0[39], keyIn_0_75, KeyWire_0[75]);
  not KeyNOTGate_0_39(G581, KeyNOTWire_0[39]);
  nand NAND2_156(G582,G462,G540);
  nand NAND2_157(KeyWire_0[76], G465,G540);
  xnor KeyGate_0_76(G583, keyIn_0_76, KeyWire_0[76]);
  nand NAND2_158(G584,G468,G543);
  nand NAND2_159(KeyWire_0[77], G471,G543);
  xnor KeyGate_0_77(KeyNOTWire_0[40], keyIn_0_77, KeyWire_0[77]);
  not KeyNOTGate_0_40(G585, KeyNOTWire_0[40]);
  nand NAND2_160(G586,G474,G546);
  nand NAND2_161(KeyWire_0[78], G477,G546);
  xnor KeyGate_0_78(G587, keyIn_0_78, KeyWire_0[78]);
  nand NAND2_162(G588,G480,G549);
  nand NAND2_163(G589,G483,G549);
  nand NAND2_164(G590,G486,G552);
  nand NAND2_165(G591,G489,G552);
  nand NAND2_166(G592,G492,G555);
  nand NAND2_167(G593,G495,G555);
  nand NAND2_168(G594,G498,G558);
  nand NAND2_169(G595,G501,G558);
  nand NAND2_170(KeyWire_0[79], G504,G561);
  xnor KeyGate_0_79(G596, keyIn_0_79, KeyWire_0[79]);
  nand NAND2_171(KeyWire_0[80], G507,G561);
  xnor KeyGate_0_80(KeyNOTWire_0[41], keyIn_0_80, KeyWire_0[80]);
  not KeyNOTGate_0_41(G597, KeyNOTWire_0[41]);
  nand NAND2_172(G598,G510,G564);
  nand NAND2_173(KeyWire_0[81], G513,G564);
  xnor KeyGate_0_81(KeyNOTWire_0[42], keyIn_0_81, KeyWire_0[81]);
  not KeyNOTGate_0_42(G599, KeyNOTWire_0[42]);
  nand NAND2_174(KeyWire_0[82], G516,G567);
  xnor KeyGate_0_82(KeyNOTWire_0[43], keyIn_0_82, KeyWire_0[82]);
  not KeyNOTGate_0_43(G600, KeyNOTWire_0[43]);
  nand NAND2_175(G601,G519,G567);
  nand NAND2_176(KeyWire_0[83], G570,G571);
  xor KeyGate_0_83(G602, keyIn_0_83, KeyWire_0[83]);
  nand NAND2_177(KeyWire_0[84], G572,G573);
  xor KeyGate_0_84(G607, keyIn_0_84, KeyWire_0[84]);
  nand NAND2_178(KeyWire_0[85], G574,G575);
  xor KeyGate_0_85(G612, keyIn_0_85, KeyWire_0[85]);
  nand NAND2_179(KeyWire_0[86], G576,G577);
  xor KeyGate_0_86(KeyNOTWire_0[44], keyIn_0_86, KeyWire_0[86]);
  not KeyNOTGate_0_44(G617, KeyNOTWire_0[44]);
  nand NAND2_180(KeyWire_0[87], G578,G579);
  xor KeyGate_0_87(KeyNOTWire_0[45], keyIn_0_87, KeyWire_0[87]);
  not KeyNOTGate_0_45(G622, KeyNOTWire_0[45]);
  nand NAND2_181(KeyWire_0[88], G580,G581);
  xnor KeyGate_0_88(G627, keyIn_0_88, KeyWire_0[88]);
  nand NAND2_182(G632,G582,G583);
  nand NAND2_183(KeyWire_0[89], G584,G585);
  xnor KeyGate_0_89(G637, keyIn_0_89, KeyWire_0[89]);
  nand NAND2_184(G642,G586,G587);
  nand NAND2_185(KeyWire_0[90], G588,G589);
  xnor KeyGate_0_90(KeyNOTWire_0[46], keyIn_0_90, KeyWire_0[90]);
  not KeyNOTGate_0_46(G645, KeyNOTWire_0[46]);
  nand NAND2_186(KeyWire_0[91], G590,G591);
  xor KeyGate_0_91(KeyNOTWire_0[47], keyIn_0_91, KeyWire_0[91]);
  not KeyNOTGate_0_47(G648, KeyNOTWire_0[47]);
  nand NAND2_187(G651,G592,G593);
  nand NAND2_188(KeyWire_0[92], G594,G595);
  xor KeyGate_0_92(G654, keyIn_0_92, KeyWire_0[92]);
  nand NAND2_189(KeyWire_0[93], G596,G597);
  xnor KeyGate_0_93(G657, keyIn_0_93, KeyWire_0[93]);
  nand NAND2_190(KeyWire_0[94], G598,G599);
  xor KeyGate_0_94(G660, keyIn_0_94, KeyWire_0[94]);
  nand NAND2_191(KeyWire_0[95], G600,G601);
  xnor KeyGate_0_95(G663, keyIn_0_95, KeyWire_0[95]);
  nand NAND2_192(G666,G602,G607);
  nand NAND2_193(KeyWire_0[96], G612,G617);
  xnor KeyGate_0_96(KeyNOTWire_0[48], keyIn_0_96, KeyWire_0[96]);
  not KeyNOTGate_0_48(G669, KeyNOTWire_0[48]);
  nand NAND2_194(G672,G602,G612);
  nand NAND2_195(G675,G607,G617);
  nand NAND2_196(G678,G622,G627);
  nand NAND2_197(G681,G632,G637);
  nand NAND2_198(KeyWire_0[97], G622,G632);
  xor KeyGate_0_97(G684, keyIn_0_97, KeyWire_0[97]);
  nand NAND2_199(KeyWire_0[98], G627,G637);
  xnor KeyGate_0_98(KeyNOTWire_0[49], keyIn_0_98, KeyWire_0[98]);
  not KeyNOTGate_0_49(G687, KeyNOTWire_0[49]);
  nand NAND2_200(KeyWire_0[99], G602,G666);
  xnor KeyGate_0_99(G690, keyIn_0_99, KeyWire_0[99]);
  nand NAND2_201(G691,G607,G666);
  nand NAND2_202(G692,G612,G669);
  nand NAND2_203(KeyWire_0[100], G617,G669);
  xor KeyGate_0_100(KeyNOTWire_0[50], keyIn_0_100, KeyWire_0[100]);
  not KeyNOTGate_0_50(G693, KeyNOTWire_0[50]);
  nand NAND2_204(G694,G602,G672);
  nand NAND2_205(G695,G612,G672);
  nand NAND2_206(G696,G607,G675);
  nand NAND2_207(KeyWire_0[101], G617,G675);
  xnor KeyGate_0_101(KeyNOTWire_0[51], keyIn_0_101, KeyWire_0[101]);
  not KeyNOTGate_0_51(G697, KeyNOTWire_0[51]);
  nand NAND2_208(KeyWire_0[102], G622,G678);
  xnor KeyGate_0_102(KeyNOTWire_0[52], keyIn_0_102, KeyWire_0[102]);
  not KeyNOTGate_0_52(G698, KeyNOTWire_0[52]);
  nand NAND2_209(KeyWire_0[103], G627,G678);
  xor KeyGate_0_103(KeyNOTWire_0[53], keyIn_0_103, KeyWire_0[103]);
  not KeyNOTGate_0_53(G699, KeyNOTWire_0[53]);
  nand NAND2_210(KeyWire_0[104], G632,G681);
  xor KeyGate_0_104(G700, keyIn_0_104, KeyWire_0[104]);
  nand NAND2_211(KeyWire_0[105], G637,G681);
  xnor KeyGate_0_105(G701, keyIn_0_105, KeyWire_0[105]);
  nand NAND2_212(G702,G622,G684);
  nand NAND2_213(G703,G632,G684);
  nand NAND2_214(KeyWire_0[106], G627,G687);
  xor KeyGate_0_106(G704, keyIn_0_106, KeyWire_0[106]);
  nand NAND2_215(G705,G637,G687);
  nand NAND2_216(G706,G690,G691);
  nand NAND2_217(KeyWire_0[107], G692,G693);
  xor KeyGate_0_107(KeyNOTWire_0[54], keyIn_0_107, KeyWire_0[107]);
  not KeyNOTGate_0_54(G709, KeyNOTWire_0[54]);
  nand NAND2_218(KeyWire_0[108], G694,G695);
  xnor KeyGate_0_108(KeyNOTWire_0[55], keyIn_0_108, KeyWire_0[108]);
  not KeyNOTGate_0_55(G712, KeyNOTWire_0[55]);
  nand NAND2_219(KeyWire_0[109], G696,G697);
  xnor KeyGate_0_109(G715, keyIn_0_109, KeyWire_0[109]);
  nand NAND2_220(KeyWire_0[110], G698,G699);
  xor KeyGate_0_110(KeyNOTWire_0[56], keyIn_0_110, KeyWire_0[110]);
  not KeyNOTGate_0_56(G718, KeyNOTWire_0[56]);
  nand NAND2_221(KeyWire_0[111], G700,G701);
  xnor KeyGate_0_111(G721, keyIn_0_111, KeyWire_0[111]);
  nand NAND2_222(G724,G702,G703);
  nand NAND2_223(G727,G704,G705);
  nand NAND2_224(G730,G242,G718);
  nand NAND2_225(G733,G245,G721);
  nand NAND2_226(G736,G248,G724);
  nand NAND2_227(KeyWire_0[112], G251,G727);
  xor KeyGate_0_112(KeyNOTWire_0[57], keyIn_0_112, KeyWire_0[112]);
  not KeyNOTGate_0_57(G739, KeyNOTWire_0[57]);
  nand NAND2_228(G742,G254,G706);
  nand NAND2_229(KeyWire_0[113], G257,G709);
  xor KeyGate_0_113(KeyNOTWire_0[58], keyIn_0_113, KeyWire_0[113]);
  not KeyNOTGate_0_58(G745, KeyNOTWire_0[58]);
  nand NAND2_230(KeyWire_0[114], G260,G712);
  xor KeyGate_0_114(KeyNOTWire_0[59], keyIn_0_114, KeyWire_0[114]);
  not KeyNOTGate_0_59(G748, KeyNOTWire_0[59]);
  nand NAND2_231(G751,G263,G715);
  nand NAND2_232(KeyWire_0[115], G242,G730);
  xnor KeyGate_0_115(KeyNOTWire_0[60], keyIn_0_115, KeyWire_0[115]);
  not KeyNOTGate_0_60(G754, KeyNOTWire_0[60]);
  nand NAND2_233(KeyWire_0[116], G718,G730);
  xor KeyGate_0_116(KeyNOTWire_0[61], keyIn_0_116, KeyWire_0[116]);
  not KeyNOTGate_0_61(G755, KeyNOTWire_0[61]);
  nand NAND2_234(G756,G245,G733);
  nand NAND2_235(G757,G721,G733);
  nand NAND2_236(G758,G248,G736);
  nand NAND2_237(G759,G724,G736);
  nand NAND2_238(G760,G251,G739);
  nand NAND2_239(KeyWire_0[117], G727,G739);
  xnor KeyGate_0_117(G761, keyIn_0_117, KeyWire_0[117]);
  nand NAND2_240(G762,G254,G742);
  nand NAND2_241(KeyWire_0[118], G706,G742);
  xor KeyGate_0_118(KeyNOTWire_0[62], keyIn_0_118, KeyWire_0[118]);
  not KeyNOTGate_0_62(G763, KeyNOTWire_0[62]);
  nand NAND2_242(KeyWire_0[119], G257,G745);
  xor KeyGate_0_119(G764, keyIn_0_119, KeyWire_0[119]);
  nand NAND2_243(KeyWire_0[120], G709,G745);
  xnor KeyGate_0_120(KeyNOTWire_0[63], keyIn_0_120, KeyWire_0[120]);
  not KeyNOTGate_0_63(G765, KeyNOTWire_0[63]);
  nand NAND2_244(KeyWire_0[121], G260,G748);
  xnor KeyGate_0_121(G766, keyIn_0_121, KeyWire_0[121]);
  nand NAND2_245(G767,G712,G748);
  nand NAND2_246(G768,G263,G751);
  nand NAND2_247(KeyWire_0[122], G715,G751);
  xor KeyGate_0_122(G769, keyIn_0_122, KeyWire_0[122]);
  nand NAND2_248(KeyWire_0[123], G754,G755);
  xnor KeyGate_0_123(KeyNOTWire_0[64], keyIn_0_123, KeyWire_0[123]);
  not KeyNOTGate_0_64(G770, KeyNOTWire_0[64]);
  nand NAND2_249(KeyWire_0[124], G756,G757);
  xnor KeyGate_0_124(KeyNOTWire_0[65], keyIn_0_124, KeyWire_0[124]);
  not KeyNOTGate_0_65(G773, KeyNOTWire_0[65]);
  nand NAND2_250(G776,G758,G759);
  nand NAND2_251(KeyWire_0[125], G760,G761);
  xnor KeyGate_0_125(KeyNOTWire_0[66], keyIn_0_125, KeyWire_0[125]);
  not KeyNOTGate_0_66(G779, KeyNOTWire_0[66]);
  nand NAND2_252(G782,G762,G763);
  nand NAND2_253(G785,G764,G765);
  nand NAND2_254(G788,G766,G767);
  nand NAND2_255(KeyWire_0[126], G768,G769);
  xnor KeyGate_0_126(KeyNOTWire_0[67], keyIn_0_126, KeyWire_0[126]);
  not KeyNOTGate_0_67(G791, KeyNOTWire_0[67]);
  nand NAND2_256(KeyWire_0[127], G642,G770);
  xor KeyGate_0_127(G794, keyIn_0_127, KeyWire_0[127]);
  nand NAND2_257(KeyWire_0[128], G645,G773);
  xnor KeyGate_0_128(G797, keyIn_0_128, KeyWire_0[128]);
  nand NAND2_258(G800,G648,G776);
  nand NAND2_259(G803,G651,G779);
  nand NAND2_260(KeyWire_0[129], G654,G782);
  xnor KeyGate_0_129(G806, keyIn_0_129, KeyWire_0[129]);
  nand NAND2_261(KeyWire_0[130], G657,G785);
  xor KeyGate_0_130(KeyNOTWire_0[68], keyIn_0_130, KeyWire_0[130]);
  not KeyNOTGate_0_68(G809, KeyNOTWire_0[68]);
  nand NAND2_262(G812,G660,G788);
  nand NAND2_263(G815,G663,G791);
  nand NAND2_264(KeyWire_0[131], G642,G794);
  xor KeyGate_0_131(KeyNOTWire_0[69], keyIn_0_131, KeyWire_0[131]);
  not KeyNOTGate_0_69(G818, KeyNOTWire_0[69]);
  nand NAND2_265(G819,G770,G794);
  nand NAND2_266(KeyWire_0[132], G645,G797);
  xnor KeyGate_0_132(KeyNOTWire_0[70], keyIn_0_132, KeyWire_0[132]);
  not KeyNOTGate_0_70(G820, KeyNOTWire_0[70]);
  nand NAND2_267(G821,G773,G797);
  nand NAND2_268(KeyWire_0[133], G648,G800);
  xor KeyGate_0_133(KeyNOTWire_0[71], keyIn_0_133, KeyWire_0[133]);
  not KeyNOTGate_0_71(G822, KeyNOTWire_0[71]);
  nand NAND2_269(KeyWire_0[134], G776,G800);
  xnor KeyGate_0_134(KeyNOTWire_0[72], keyIn_0_134, KeyWire_0[134]);
  not KeyNOTGate_0_72(G823, KeyNOTWire_0[72]);
  nand NAND2_270(G824,G651,G803);
  nand NAND2_271(KeyWire_0[135], G779,G803);
  xnor KeyGate_0_135(KeyNOTWire_0[73], keyIn_0_135, KeyWire_0[135]);
  not KeyNOTGate_0_73(G825, KeyNOTWire_0[73]);
  nand NAND2_272(G826,G654,G806);
  nand NAND2_273(KeyWire_0[136], G782,G806);
  xor KeyGate_0_136(KeyNOTWire_0[74], keyIn_0_136, KeyWire_0[136]);
  not KeyNOTGate_0_74(G827, KeyNOTWire_0[74]);
  nand NAND2_274(G828,G657,G809);
  nand NAND2_275(KeyWire_0[137], G785,G809);
  xnor KeyGate_0_137(KeyNOTWire_0[75], keyIn_0_137, KeyWire_0[137]);
  not KeyNOTGate_0_75(G829, KeyNOTWire_0[75]);
  nand NAND2_276(G830,G660,G812);
  nand NAND2_277(G831,G788,G812);
  nand NAND2_278(G832,G663,G815);
  nand NAND2_279(G833,G791,G815);
  nand NAND2_280(G834,G818,G819);
  nand NAND2_281(KeyWire_0[138], G820,G821);
  xnor KeyGate_0_138(KeyNOTWire_0[76], keyIn_0_138, KeyWire_0[138]);
  not KeyNOTGate_0_76(G847, KeyNOTWire_0[76]);
  nand NAND2_282(KeyWire_0[139], G822,G823);
  xnor KeyGate_0_139(G860, keyIn_0_139, KeyWire_0[139]);
  nand NAND2_283(KeyWire_0[140], G824,G825);
  xor KeyGate_0_140(G873, keyIn_0_140, KeyWire_0[140]);
  nand NAND2_284(KeyWire_0[141], G828,G829);
  xnor KeyGate_0_141(G886, keyIn_0_141, KeyWire_0[141]);
  nand NAND2_285(KeyWire_0[142], G832,G833);
  xor KeyGate_0_142(G899, keyIn_0_142, KeyWire_0[142]);
  nand NAND2_286(G912,G830,G831);
  nand NAND2_287(G925,G826,G827);
  not NOT_0(KeyWire_0[143], G834);
  xor KeyGate_0_143(KeyNOTWire_0[77], keyIn_0_143, KeyWire_0[143]);
  not KeyNOTGate_0_77(G938, KeyNOTWire_0[77]);
  not NOT_1(G939,G847);
  not NOT_2(KeyWire_0[144], G860);
  xor KeyGate_0_144(G940, keyIn_0_144, KeyWire_0[144]);
  not NOT_3(G941,G834);
  not NOT_4(G942,G847);
  not NOT_5(G943,G873);
  not NOT_6(KeyWire_0[145], G834);
  xnor KeyGate_0_145(KeyNOTWire_0[78], keyIn_0_145, KeyWire_0[145]);
  not KeyNOTGate_0_78(G944, KeyNOTWire_0[78]);
  not NOT_7(G945,G860);
  not NOT_8(KeyWire_0[146], G873);
  xnor KeyGate_0_146(KeyNOTWire_0[79], keyIn_0_146, KeyWire_0[146]);
  not KeyNOTGate_0_79(G946, KeyNOTWire_0[79]);
  not NOT_9(KeyWire_0[147], G847);
  xnor KeyGate_0_147(G947, keyIn_0_147, KeyWire_0[147]);
  not NOT_10(KeyWire_0[148], G860);
  xnor KeyGate_0_148(KeyNOTWire_0[80], keyIn_0_148, KeyWire_0[148]);
  not KeyNOTGate_0_80(G948, KeyNOTWire_0[80]);
  not NOT_11(G949,G873);
  not NOT_12(G950,G886);
  not NOT_13(G951,G899);
  not NOT_14(KeyWire_0[149], G886);
  xor KeyGate_0_149(KeyNOTWire_0[81], keyIn_0_149, KeyWire_0[149]);
  not KeyNOTGate_0_81(G952, KeyNOTWire_0[81]);
  not NOT_15(G953,G912);
  not NOT_16(G954,G925);
  not NOT_17(KeyWire_0[150], G899);
  xnor KeyGate_0_150(G955, keyIn_0_150, KeyWire_0[150]);
  not NOT_18(G956,G925);
  not NOT_19(G957,G912);
  not NOT_20(KeyWire_0[151], G925);
  xor KeyGate_0_151(G958, keyIn_0_151, KeyWire_0[151]);
  not NOT_21(KeyWire_0[152], G886);
  xnor KeyGate_0_152(G959, keyIn_0_152, KeyWire_0[152]);
  not NOT_22(G960,G912);
  not NOT_23(G961,G925);
  not NOT_24(G962,G886);
  not NOT_25(G963,G899);
  not NOT_26(KeyWire_0[153], G925);
  xor KeyGate_0_153(G964, keyIn_0_153, KeyWire_0[153]);
  not NOT_27(G965,G912);
  not NOT_28(KeyWire_0[154], G899);
  xnor KeyGate_0_154(G966, keyIn_0_154, KeyWire_0[154]);
  not NOT_29(KeyWire_0[155], G886);
  xor KeyGate_0_155(KeyNOTWire_0[82], keyIn_0_155, KeyWire_0[155]);
  not KeyNOTGate_0_82(G967, KeyNOTWire_0[82]);
  not NOT_30(KeyWire_0[156], G912);
  xnor KeyGate_0_156(KeyNOTWire_0[83], keyIn_0_156, KeyWire_0[156]);
  not KeyNOTGate_0_83(G968, KeyNOTWire_0[83]);
  not NOT_31(G969,G899);
  not NOT_32(G970,G847);
  not NOT_33(G971,G873);
  not NOT_34(G972,G847);
  not NOT_35(G973,G860);
  not NOT_36(KeyWire_0[157], G834);
  xnor KeyGate_0_157(KeyNOTWire_0[84], keyIn_0_157, KeyWire_0[157]);
  not KeyNOTGate_0_84(G974, KeyNOTWire_0[84]);
  not NOT_37(G975,G873);
  not NOT_38(G976,G834);
  not NOT_39(G977,G860);
  and AND4_0(G978,G938,G939,G940,G873);
  and AND4_1(KeyWire_0[158], G941,G942,G860,G943);
  xor KeyGate_0_158(KeyNOTWire_0[85], keyIn_0_158, KeyWire_0[158]);
  not KeyNOTGate_0_85(G979, KeyNOTWire_0[85]);
  and AND4_2(G980,G944,G847,G945,G946);
  and AND4_3(KeyWire_0[159], G834,G947,G948,G949);
  xnor KeyGate_0_159(KeyNOTWire_0[86], keyIn_0_159, KeyWire_0[159]);
  not KeyNOTGate_0_86(G981, KeyNOTWire_0[86]);
  and AND4_4(KeyWire_0[160], G958,G959,G960,G899);
  xnor KeyGate_0_160(G982, keyIn_0_160, KeyWire_0[160]);
  and AND4_5(KeyWire_0[161], G961,G962,G912,G963);
  xor KeyGate_0_161(G983, keyIn_0_161, KeyWire_0[161]);
  and AND4_6(KeyWire_0[162], G964,G886,G965,G966);
  xnor KeyGate_0_162(G984, keyIn_0_162, KeyWire_0[162]);
  and AND4_7(KeyWire_0[163], G925,G967,G968,G969);
  xnor KeyGate_0_163(G985, keyIn_0_163, KeyWire_0[163]);
  or OR4_0(KeyWire_0[164], G978,G979,G980,G981);
  xor KeyGate_0_164(G986, keyIn_0_164, KeyWire_0[164]);
  or OR4_1(G991,G982,G983,G984,G985);
  and AND5_0(KeyWire_0[165], G925,G950,G912,G951,G986);
  xor KeyGate_0_165(KeyNOTWire_0[87], keyIn_0_165, KeyWire_0[165]);
  not KeyNOTGate_0_87(G996, KeyNOTWire_0[87]);
  and AND5_1(G1001,G925,G952,G953,G899,G986);
  and AND5_2(KeyWire_0[166], G954,G886,G912,G955,G986);
  xnor KeyGate_0_166(KeyNOTWire_0[88], keyIn_0_166, KeyWire_0[166]);
  not KeyNOTGate_0_88(G1006, KeyNOTWire_0[88]);
  and AND5_3(KeyWire_0[167], G956,G886,G957,G899,G986);
  xnor KeyGate_0_167(G1011, keyIn_0_167, KeyWire_0[167]);
  and AND5_4(G1016,G834,G970,G860,G971,G991);
  and AND5_5(KeyWire_0[168], G834,G972,G973,G873,G991);
  xor KeyGate_0_168(G1021, keyIn_0_168, KeyWire_0[168]);
  and AND5_6(G1026,G974,G847,G860,G975,G991);
  and AND5_7(KeyWire_0[169], G976,G847,G977,G873,G991);
  xnor KeyGate_0_169(G1031, keyIn_0_169, KeyWire_0[169]);
  and AND2_8(G1036,G834,G996);
  and AND2_9(KeyWire_0[170], G847,G996);
  xnor KeyGate_0_170(KeyNOTWire_0[89], keyIn_0_170, KeyWire_0[170]);
  not KeyNOTGate_0_89(G1039, KeyNOTWire_0[89]);
  and AND2_10(KeyWire_0[171], G860,G996);
  xnor KeyGate_0_171(G1042, keyIn_0_171, KeyWire_0[171]);
  and AND2_11(G1045,G873,G996);
  and AND2_12(KeyWire_0[172], G834,G1001);
  xnor KeyGate_0_172(KeyNOTWire_0[90], keyIn_0_172, KeyWire_0[172]);
  not KeyNOTGate_0_90(G1048, KeyNOTWire_0[90]);
  and AND2_13(KeyWire_0[173], G847,G1001);
  xor KeyGate_0_173(KeyNOTWire_0[91], keyIn_0_173, KeyWire_0[173]);
  not KeyNOTGate_0_91(G1051, KeyNOTWire_0[91]);
  and AND2_14(G1054,G860,G1001);
  and AND2_15(KeyWire_0[174], G873,G1001);
  xor KeyGate_0_174(KeyNOTWire_0[92], keyIn_0_174, KeyWire_0[174]);
  not KeyNOTGate_0_92(G1057, KeyNOTWire_0[92]);
  and AND2_16(G1060,G834,G1006);
  and AND2_17(G1063,G847,G1006);
  and AND2_18(G1066,G860,G1006);
  and AND2_19(G1069,G873,G1006);
  and AND2_20(G1072,G834,G1011);
  and AND2_21(G1075,G847,G1011);
  and AND2_22(G1078,G860,G1011);
  and AND2_23(G1081,G873,G1011);
  and AND2_24(KeyWire_0[175], G925,G1016);
  xor KeyGate_0_175(KeyNOTWire_0[93], keyIn_0_175, KeyWire_0[175]);
  not KeyNOTGate_0_93(G1084, KeyNOTWire_0[93]);
  and AND2_25(KeyWire_0[176], G886,G1016);
  xnor KeyGate_0_176(G1087, keyIn_0_176, KeyWire_0[176]);
  and AND2_26(G1090,G912,G1016);
  and AND2_27(G1093,G899,G1016);
  and AND2_28(KeyWire_0[177], G925,G1021);
  xnor KeyGate_0_177(KeyNOTWire_0[94], keyIn_0_177, KeyWire_0[177]);
  not KeyNOTGate_0_94(G1096, KeyNOTWire_0[94]);
  and AND2_29(G1099,G886,G1021);
  and AND2_30(G1102,G912,G1021);
  and AND2_31(KeyWire_0[178], G899,G1021);
  xnor KeyGate_0_178(KeyNOTWire_0[95], keyIn_0_178, KeyWire_0[178]);
  not KeyNOTGate_0_95(G1105, KeyNOTWire_0[95]);
  and AND2_32(KeyWire_0[179], G925,G1026);
  xor KeyGate_0_179(KeyNOTWire_0[96], keyIn_0_179, KeyWire_0[179]);
  not KeyNOTGate_0_96(G1108, KeyNOTWire_0[96]);
  and AND2_33(G1111,G886,G1026);
  and AND2_34(G1114,G912,G1026);
  and AND2_35(G1117,G899,G1026);
  and AND2_36(G1120,G925,G1031);
  and AND2_37(G1123,G886,G1031);
  and AND2_38(KeyWire_0[180], G912,G1031);
  xor KeyGate_0_180(G1126, keyIn_0_180, KeyWire_0[180]);
  and AND2_39(KeyWire_0[181], G899,G1031);
  xor KeyGate_0_181(KeyNOTWire_0[97], keyIn_0_181, KeyWire_0[181]);
  not KeyNOTGate_0_97(G1129, KeyNOTWire_0[97]);
  nand NAND2_288(G1132,G1,G1036);
  nand NAND2_289(KeyWire_0[182], G2,G1039);
  xnor KeyGate_0_182(KeyNOTWire_0[98], keyIn_0_182, KeyWire_0[182]);
  not KeyNOTGate_0_98(G1135, KeyNOTWire_0[98]);
  nand NAND2_290(G1138,G3,G1042);
  nand NAND2_291(G1141,G4,G1045);
  nand NAND2_292(G1144,G5,G1048);
  nand NAND2_293(KeyWire_0[183], G6,G1051);
  xnor KeyGate_0_183(G1147, keyIn_0_183, KeyWire_0[183]);
  nand NAND2_294(KeyWire_0[184], G7,G1054);
  xnor KeyGate_0_184(G1150, keyIn_0_184, KeyWire_0[184]);
  nand NAND2_295(KeyWire_0[185], G8,G1057);
  xnor KeyGate_0_185(G1153, keyIn_0_185, KeyWire_0[185]);
  nand NAND2_296(KeyWire_0[186], G9,G1060);
  xor KeyGate_0_186(KeyNOTWire_0[99], keyIn_0_186, KeyWire_0[186]);
  not KeyNOTGate_0_99(G1156, KeyNOTWire_0[99]);
  nand NAND2_297(KeyWire_0[187], G10,G1063);
  xnor KeyGate_0_187(KeyNOTWire_0[100], keyIn_0_187, KeyWire_0[187]);
  not KeyNOTGate_0_100(G1159, KeyNOTWire_0[100]);
  nand NAND2_298(G1162,G11,G1066);
  nand NAND2_299(KeyWire_0[188], G12,G1069);
  xnor KeyGate_0_188(G1165, keyIn_0_188, KeyWire_0[188]);
  nand NAND2_300(KeyWire_0[189], G13,G1072);
  xor KeyGate_0_189(KeyNOTWire_0[101], keyIn_0_189, KeyWire_0[189]);
  not KeyNOTGate_0_101(G1168, KeyNOTWire_0[101]);
  nand NAND2_301(KeyWire_0[190], G14,G1075);
  xor KeyGate_0_190(G1171, keyIn_0_190, KeyWire_0[190]);
  nand NAND2_302(KeyWire_0[191], G15,G1078);
  xnor KeyGate_0_191(G1174, keyIn_0_191, KeyWire_0[191]);
  nand NAND2_303(KeyWire_0[192], G16,G1081);
  xor KeyGate_0_192(KeyNOTWire_0[102], keyIn_0_192, KeyWire_0[192]);
  not KeyNOTGate_0_102(G1177, KeyNOTWire_0[102]);
  nand NAND2_304(G1180,G17,G1084);
  nand NAND2_305(KeyWire_0[193], G18,G1087);
  xnor KeyGate_0_193(KeyNOTWire_0[103], keyIn_0_193, KeyWire_0[193]);
  not KeyNOTGate_0_103(G1183, KeyNOTWire_0[103]);
  nand NAND2_306(KeyWire_0[194], G19,G1090);
  xor KeyGate_0_194(G1186, keyIn_0_194, KeyWire_0[194]);
  nand NAND2_307(G1189,G20,G1093);
  nand NAND2_308(KeyWire_0[195], G21,G1096);
  xor KeyGate_0_195(KeyNOTWire_0[104], keyIn_0_195, KeyWire_0[195]);
  not KeyNOTGate_0_104(G1192, KeyNOTWire_0[104]);
  nand NAND2_309(G1195,G22,G1099);
  nand NAND2_310(KeyWire_0[196], G23,G1102);
  xor KeyGate_0_196(KeyNOTWire_0[105], keyIn_0_196, KeyWire_0[196]);
  not KeyNOTGate_0_105(G1198, KeyNOTWire_0[105]);
  nand NAND2_311(KeyWire_0[197], G24,G1105);
  xnor KeyGate_0_197(KeyNOTWire_0[106], keyIn_0_197, KeyWire_0[197]);
  not KeyNOTGate_0_106(G1201, KeyNOTWire_0[106]);
  nand NAND2_312(KeyWire_0[198], G25,G1108);
  xor KeyGate_0_198(KeyNOTWire_0[107], keyIn_0_198, KeyWire_0[198]);
  not KeyNOTGate_0_107(G1204, KeyNOTWire_0[107]);
  nand NAND2_313(G1207,G26,G1111);
  nand NAND2_314(G1210,G27,G1114);
  nand NAND2_315(G1213,G28,G1117);
  nand NAND2_316(KeyWire_0[199], G29,G1120);
  xor KeyGate_0_199(KeyNOTWire_0[108], keyIn_0_199, KeyWire_0[199]);
  not KeyNOTGate_0_108(G1216, KeyNOTWire_0[108]);
  nand NAND2_317(G1219,G30,G1123);
  nand NAND2_318(KeyWire_0[200], G31,G1126);
  xnor KeyGate_0_200(G1222, keyIn_0_200, KeyWire_0[200]);
  nand NAND2_319(KeyWire_0[201], G32,G1129);
  xor KeyGate_0_201(G1225, keyIn_0_201, KeyWire_0[201]);
  nand NAND2_320(KeyWire_0[202], G1,G1132);
  xnor KeyGate_0_202(G1228, keyIn_0_202, KeyWire_0[202]);
  nand NAND2_321(KeyWire_0[203], G1036,G1132);
  xnor KeyGate_0_203(G1229, keyIn_0_203, KeyWire_0[203]);
  nand NAND2_322(G1230,G2,G1135);
  nand NAND2_323(G1231,G1039,G1135);
  nand NAND2_324(G1232,G3,G1138);
  nand NAND2_325(G1233,G1042,G1138);
  nand NAND2_326(G1234,G4,G1141);
  nand NAND2_327(G1235,G1045,G1141);
  nand NAND2_328(G1236,G5,G1144);
  nand NAND2_329(G1237,G1048,G1144);
  nand NAND2_330(G1238,G6,G1147);
  nand NAND2_331(G1239,G1051,G1147);
  nand NAND2_332(G1240,G7,G1150);
  nand NAND2_333(KeyWire_0[204], G1054,G1150);
  xor KeyGate_0_204(G1241, keyIn_0_204, KeyWire_0[204]);
  nand NAND2_334(G1242,G8,G1153);
  nand NAND2_335(KeyWire_0[205], G1057,G1153);
  xor KeyGate_0_205(KeyNOTWire_0[109], keyIn_0_205, KeyWire_0[205]);
  not KeyNOTGate_0_109(G1243, KeyNOTWire_0[109]);
  nand NAND2_336(KeyWire_0[206], G9,G1156);
  xor KeyGate_0_206(KeyNOTWire_0[110], keyIn_0_206, KeyWire_0[206]);
  not KeyNOTGate_0_110(G1244, KeyNOTWire_0[110]);
  nand NAND2_337(G1245,G1060,G1156);
  nand NAND2_338(G1246,G10,G1159);
  nand NAND2_339(KeyWire_0[207], G1063,G1159);
  xnor KeyGate_0_207(G1247, keyIn_0_207, KeyWire_0[207]);
  nand NAND2_340(G1248,G11,G1162);
  nand NAND2_341(G1249,G1066,G1162);
  nand NAND2_342(G1250,G12,G1165);
  nand NAND2_343(G1251,G1069,G1165);
  nand NAND2_344(G1252,G13,G1168);
  nand NAND2_345(KeyWire_0[208], G1072,G1168);
  xnor KeyGate_0_208(G1253, keyIn_0_208, KeyWire_0[208]);
  nand NAND2_346(G1254,G14,G1171);
  nand NAND2_347(KeyWire_0[209], G1075,G1171);
  xor KeyGate_0_209(G1255, keyIn_0_209, KeyWire_0[209]);
  nand NAND2_348(KeyWire_0[210], G15,G1174);
  xnor KeyGate_0_210(KeyNOTWire_0[111], keyIn_0_210, KeyWire_0[210]);
  not KeyNOTGate_0_111(G1256, KeyNOTWire_0[111]);
  nand NAND2_349(KeyWire_0[211], G1078,G1174);
  xnor KeyGate_0_211(G1257, keyIn_0_211, KeyWire_0[211]);
  nand NAND2_350(G1258,G16,G1177);
  nand NAND2_351(G1259,G1081,G1177);
  nand NAND2_352(KeyWire_0[212], G17,G1180);
  xnor KeyGate_0_212(KeyNOTWire_0[112], keyIn_0_212, KeyWire_0[212]);
  not KeyNOTGate_0_112(G1260, KeyNOTWire_0[112]);
  nand NAND2_353(G1261,G1084,G1180);
  nand NAND2_354(KeyWire_0[213], G18,G1183);
  xnor KeyGate_0_213(KeyNOTWire_0[113], keyIn_0_213, KeyWire_0[213]);
  not KeyNOTGate_0_113(G1262, KeyNOTWire_0[113]);
  nand NAND2_355(G1263,G1087,G1183);
  nand NAND2_356(G1264,G19,G1186);
  nand NAND2_357(G1265,G1090,G1186);
  nand NAND2_358(KeyWire_0[214], G20,G1189);
  xor KeyGate_0_214(G1266, keyIn_0_214, KeyWire_0[214]);
  nand NAND2_359(KeyWire_0[215], G1093,G1189);
  xnor KeyGate_0_215(G1267, keyIn_0_215, KeyWire_0[215]);
  nand NAND2_360(G1268,G21,G1192);
  nand NAND2_361(G1269,G1096,G1192);
  nand NAND2_362(G1270,G22,G1195);
  nand NAND2_363(KeyWire_0[216], G1099,G1195);
  xnor KeyGate_0_216(G1271, keyIn_0_216, KeyWire_0[216]);
  nand NAND2_364(KeyWire_0[217], G23,G1198);
  xor KeyGate_0_217(KeyNOTWire_0[114], keyIn_0_217, KeyWire_0[217]);
  not KeyNOTGate_0_114(G1272, KeyNOTWire_0[114]);
  nand NAND2_365(G1273,G1102,G1198);
  nand NAND2_366(G1274,G24,G1201);
  nand NAND2_367(G1275,G1105,G1201);
  nand NAND2_368(G1276,G25,G1204);
  nand NAND2_369(G1277,G1108,G1204);
  nand NAND2_370(G1278,G26,G1207);
  nand NAND2_371(KeyWire_0[218], G1111,G1207);
  xor KeyGate_0_218(G1279, keyIn_0_218, KeyWire_0[218]);
  nand NAND2_372(G1280,G27,G1210);
  nand NAND2_373(KeyWire_0[219], G1114,G1210);
  xor KeyGate_0_219(KeyNOTWire_0[115], keyIn_0_219, KeyWire_0[219]);
  not KeyNOTGate_0_115(G1281, KeyNOTWire_0[115]);
  nand NAND2_374(G1282,G28,G1213);
  nand NAND2_375(KeyWire_0[220], G1117,G1213);
  xnor KeyGate_0_220(G1283, keyIn_0_220, KeyWire_0[220]);
  nand NAND2_376(G1284,G29,G1216);
  nand NAND2_377(KeyWire_0[221], G1120,G1216);
  xor KeyGate_0_221(KeyNOTWire_0[116], keyIn_0_221, KeyWire_0[221]);
  not KeyNOTGate_0_116(G1285, KeyNOTWire_0[116]);
  nand NAND2_378(KeyWire_0[222], G30,G1219);
  xor KeyGate_0_222(KeyNOTWire_0[117], keyIn_0_222, KeyWire_0[222]);
  not KeyNOTGate_0_117(G1286, KeyNOTWire_0[117]);
  nand NAND2_379(KeyWire_0[223], G1123,G1219);
  xor KeyGate_0_223(G1287, keyIn_0_223, KeyWire_0[223]);
  nand NAND2_380(G1288,G31,G1222);
  nand NAND2_381(G1289,G1126,G1222);
  nand NAND2_382(G1290,G32,G1225);
  nand NAND2_383(KeyWire_0[224], G1129,G1225);
  xnor KeyGate_0_224(G1291, keyIn_0_224, KeyWire_0[224]);
  nand NAND2_384(G1292,G1228,G1229);
  nand NAND2_385(G1293,G1230,G1231);
  nand NAND2_386(G1294,G1232,G1233);
  nand NAND2_387(G1295,G1234,G1235);
  nand NAND2_388(KeyWire_0[225], G1236,G1237);
  xor KeyGate_0_225(KeyNOTWire_0[118], keyIn_0_225, KeyWire_0[225]);
  not KeyNOTGate_0_118(G1296, KeyNOTWire_0[118]);
  nand NAND2_389(G1297,G1238,G1239);
  nand NAND2_390(G1298,G1240,G1241);
  nand NAND2_391(KeyWire_0[226], G1242,G1243);
  xor KeyGate_0_226(G1299, keyIn_0_226, KeyWire_0[226]);
  nand NAND2_392(KeyWire_0[227], G1244,G1245);
  xnor KeyGate_0_227(KeyNOTWire_0[119], keyIn_0_227, KeyWire_0[227]);
  not KeyNOTGate_0_119(G1300, KeyNOTWire_0[119]);
  nand NAND2_393(KeyWire_0[228], G1246,G1247);
  xnor KeyGate_0_228(G1301, keyIn_0_228, KeyWire_0[228]);
  nand NAND2_394(G1302,G1248,G1249);
  nand NAND2_395(G1303,G1250,G1251);
  nand NAND2_396(G1304,G1252,G1253);
  nand NAND2_397(KeyWire_0[229], G1254,G1255);
  xnor KeyGate_0_229(G1305, keyIn_0_229, KeyWire_0[229]);
  nand NAND2_398(G1306,G1256,G1257);
  nand NAND2_399(KeyWire_0[230], G1258,G1259);
  xnor KeyGate_0_230(KeyNOTWire_0[120], keyIn_0_230, KeyWire_0[230]);
  not KeyNOTGate_0_120(G1307, KeyNOTWire_0[120]);
  nand NAND2_400(G1308,G1260,G1261);
  nand NAND2_401(G1309,G1262,G1263);
  nand NAND2_402(KeyWire_0[231], G1264,G1265);
  xnor KeyGate_0_231(KeyNOTWire_0[121], keyIn_0_231, KeyWire_0[231]);
  not KeyNOTGate_0_121(G1310, KeyNOTWire_0[121]);
  nand NAND2_403(KeyWire_0[232], G1266,G1267);
  xor KeyGate_0_232(KeyNOTWire_0[122], keyIn_0_232, KeyWire_0[232]);
  not KeyNOTGate_0_122(G1311, KeyNOTWire_0[122]);
  nand NAND2_404(KeyWire_0[233], G1268,G1269);
  xor KeyGate_0_233(KeyNOTWire_0[123], keyIn_0_233, KeyWire_0[233]);
  not KeyNOTGate_0_123(G1312, KeyNOTWire_0[123]);
  nand NAND2_405(KeyWire_0[234], G1270,G1271);
  xor KeyGate_0_234(KeyNOTWire_0[124], keyIn_0_234, KeyWire_0[234]);
  not KeyNOTGate_0_124(G1313, KeyNOTWire_0[124]);
  nand NAND2_406(G1314,G1272,G1273);
  nand NAND2_407(G1315,G1274,G1275);
  nand NAND2_408(G1316,G1276,G1277);
  nand NAND2_409(G1317,G1278,G1279);
  nand NAND2_410(G1318,G1280,G1281);
  nand NAND2_411(G1319,G1282,G1283);
  nand NAND2_412(G1320,G1284,G1285);
  nand NAND2_413(G1321,G1286,G1287);
  nand NAND2_414(G1322,G1288,G1289);
  nand NAND2_415(KeyWire_0[235], G1290,G1291);
  xnor KeyGate_0_235(G1323, keyIn_0_235, KeyWire_0[235]);
  not NOT_40(G1324,G1292);
  not NOT_41(G1325,G1293);
  not NOT_42(KeyWire_0[236], G1294);
  xor KeyGate_0_236(KeyNOTWire_0[125], keyIn_0_236, KeyWire_0[236]);
  not KeyNOTGate_0_125(G1326, KeyNOTWire_0[125]);
  not NOT_43(KeyWire_0[237], G1295);
  xnor KeyGate_0_237(G1327, keyIn_0_237, KeyWire_0[237]);
  not NOT_44(KeyWire_0[238], G1296);
  xnor KeyGate_0_238(KeyNOTWire_0[126], keyIn_0_238, KeyWire_0[238]);
  not KeyNOTGate_0_126(G1328, KeyNOTWire_0[126]);
  not NOT_45(KeyWire_0[239], G1297);
  xor KeyGate_0_239(KeyNOTWire_0[127], keyIn_0_239, KeyWire_0[239]);
  not KeyNOTGate_0_127(G1329, KeyNOTWire_0[127]);
  not NOT_46(KeyWire_0[240], G1298);
  xnor KeyGate_0_240(G1330, keyIn_0_240, KeyWire_0[240]);
  not NOT_47(KeyWire_0[241], G1299);
  xnor KeyGate_0_241(KeyNOTWire_0[128], keyIn_0_241, KeyWire_0[241]);
  not KeyNOTGate_0_128(G1331, KeyNOTWire_0[128]);
  not NOT_48(KeyWire_0[242], G1300);
  xor KeyGate_0_242(KeyNOTWire_0[129], keyIn_0_242, KeyWire_0[242]);
  not KeyNOTGate_0_129(G1332, KeyNOTWire_0[129]);
  not NOT_49(KeyWire_0[243], G1301);
  xor KeyGate_0_243(KeyNOTWire_0[130], keyIn_0_243, KeyWire_0[243]);
  not KeyNOTGate_0_130(G1333, KeyNOTWire_0[130]);
  not NOT_50(G1334,G1302);
  not NOT_51(G1335,G1303);
  not NOT_52(KeyWire_0[244], G1304);
  xor KeyGate_0_244(KeyNOTWire_0[131], keyIn_0_244, KeyWire_0[244]);
  not KeyNOTGate_0_131(G1336, KeyNOTWire_0[131]);
  not NOT_53(KeyWire_0[245], G1305);
  xor KeyGate_0_245(G1337, keyIn_0_245, KeyWire_0[245]);
  not NOT_54(G1338,G1306);
  not NOT_55(KeyWire_0[246], G1307);
  xor KeyGate_0_246(KeyNOTWire_0[132], keyIn_0_246, KeyWire_0[246]);
  not KeyNOTGate_0_132(G1339, KeyNOTWire_0[132]);
  not NOT_56(KeyWire_0[247], G1308);
  xor KeyGate_0_247(G1340, keyIn_0_247, KeyWire_0[247]);
  not NOT_57(KeyWire_0[248], G1309);
  xnor KeyGate_0_248(G1341, keyIn_0_248, KeyWire_0[248]);
  not NOT_58(KeyWire_0[249], G1310);
  xor KeyGate_0_249(KeyNOTWire_0[133], keyIn_0_249, KeyWire_0[249]);
  not KeyNOTGate_0_133(G1342, KeyNOTWire_0[133]);
  not NOT_59(KeyWire_0[250], G1311);
  xnor KeyGate_0_250(KeyNOTWire_0[134], keyIn_0_250, KeyWire_0[250]);
  not KeyNOTGate_0_134(G1343, KeyNOTWire_0[134]);
  not NOT_60(G1344,G1312);
  not NOT_61(KeyWire_0[251], G1313);
  xnor KeyGate_0_251(KeyNOTWire_0[135], keyIn_0_251, KeyWire_0[251]);
  not KeyNOTGate_0_135(G1345, KeyNOTWire_0[135]);
  not NOT_62(KeyWire_0[252], G1314);
  xnor KeyGate_0_252(KeyNOTWire_0[136], keyIn_0_252, KeyWire_0[252]);
  not KeyNOTGate_0_136(G1346, KeyNOTWire_0[136]);
  not NOT_63(KeyWire_0[253], G1315);
  xnor KeyGate_0_253(G1347, keyIn_0_253, KeyWire_0[253]);
  not NOT_64(G1348,G1316);
  not NOT_65(G1349,G1317);
  not NOT_66(KeyWire_0[254], G1318);
  xor KeyGate_0_254(G1350, keyIn_0_254, KeyWire_0[254]);
  not NOT_67(KeyWire_0[255], G1319);
  xnor KeyGate_0_255(KeyNOTWire_0[137], keyIn_0_255, KeyWire_0[255]);
  not KeyNOTGate_0_137(G1351, KeyNOTWire_0[137]);
  not NOT_68(G1352,G1320);
  not NOT_69(G1353,G1321);
  not NOT_70(G1354,G1322);
  not NOT_71(G1355,G1323);

endmodule

