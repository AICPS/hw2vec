`timescale 1ns / 1ps
// Verilog
// c432
// Ninputs 36
// Noutputs 7
// NtotalGates 160
// NOT1 40
// NAND2 64
// NOR2 19
// AND9 3
// XOR2 18
// NAND4 14
// AND8 1
// NAND3 1

module top (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
                  N430,N431,N432,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
                  keyinput60, keyinput61, keyinput62, keyinput63,
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
        keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
        keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
        keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
        keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
        keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
                  keyinput134, keyinput135,
        keyinput136, keyinput137, keyinput138, keyinput139, keyinput140,
        keyinput141, keyinput142, keyinput143, keyinput144, keyinput145,
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150,
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155,
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160,
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165,
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170,
        keyinput171);

  input keyinput136, keyinput137, keyinput138, keyinput139, keyinput140;
  input keyinput141, keyinput142, keyinput143, keyinput144, keyinput145;
  input keyinput146, keyinput147, keyinput148, keyinput149, keyinput150;
  input keyinput151, keyinput152, keyinput153, keyinput154, keyinput155;
  input keyinput156, keyinput157, keyinput158, keyinput159, keyinput160;
  input keyinput161, keyinput162, keyinput163, keyinput164, keyinput165;
  input keyinput166, keyinput167, keyinput168, keyinput169, keyinput170;
  input keyinput171;


  input keyinput64, keyinput65, keyinput66, keyinput67, keyinput68;
  input keyinput69, keyinput70, keyinput71, keyinput72, keyinput73;
  input keyinput74, keyinput75, keyinput76, keyinput77, keyinput78;
  input keyinput79, keyinput80, keyinput81, keyinput82, keyinput83;
  input keyinput84, keyinput85, keyinput86, keyinput87, keyinput88;
  input keyinput89, keyinput90, keyinput91, keyinput92, keyinput93;
  input keyinput94, keyinput95, keyinput96, keyinput97, keyinput98;
  input keyinput99, keyinput100, keyinput101, keyinput102, keyinput103;
  input keyinput104, keyinput105, keyinput106, keyinput107, keyinput108;
  input keyinput109, keyinput110, keyinput111, keyinput112, keyinput113;
  input keyinput114, keyinput115, keyinput116, keyinput117, keyinput118;
  input keyinput119, keyinput120, keyinput121, keyinput122, keyinput123;
  input keyinput124, keyinput125, keyinput126, keyinput127, keyinput128;
  input keyinput129, keyinput130, keyinput131, keyinput132, keyinput133;
  input keyinput134, keyinput135;

  wire KeyWire_0_1 , KeyWire_0_2;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31, keyinput32, keyinput33, keyinput34;
  input keyinput35, keyinput36, keyinput37, keyinput38, keyinput39;
  input keyinput40, keyinput41, keyinput42, keyinput43, keyinput44;
  input keyinput45, keyinput46, keyinput47, keyinput48, keyinput49;
  input keyinput50, keyinput51, keyinput52, keyinput53, keyinput54;
  input keyinput55, keyinput56, keyinput57, keyinput58, keyinput59;
  input keyinput60, keyinput61, keyinput62, keyinput63;

  wire [0:63] keyinput_Wire_0;
  wire [0:37] KeyNOTWire_0;

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;

output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429;

  not NOT1_1 (keyinput_Wire_0[0], N1);
  xnor keyGate_0_0(KeyNOTWire_0[0], keyinput0, keyinput_Wire_0[0]);
  not KeyNOTGate_0_0(N118, KeyNOTWire_0[0]);
not NOT1_2 (N119, N4);
  not NOT1_3 (keyinput_Wire_0[1], N11);
  xnor keyGate_0_1(KeyNOTWire_0[1], keyinput1, keyinput_Wire_0[1]);
  not KeyNOTGate_0_1(N122, KeyNOTWire_0[1]);
not NOT1_4 (N123, N17);
  not NOT1_5 (keyinput_Wire_0[2], N24);
  xnor keyGate_0_2(N126, keyinput2, keyinput_Wire_0[2]);
not NOT1_6 (N127, N30);
  not NOT1_7 (keyinput_Wire_0[3], N37);
  xor keyGate_0_3(N130, keyinput3, keyinput_Wire_0[3]);
not NOT1_8 (N131, N43);
  not NOT1_9 (keyinput_Wire_0[4], N50);
  xor keyGate_0_4(KeyNOTWire_0[2], keyinput4, keyinput_Wire_0[4]);
  not KeyNOTGate_0_2(N134, KeyNOTWire_0[2]);
not NOT1_10 (N135, N56);
  not NOT1_11 (keyinput_Wire_0[5], N63);
  xor keyGate_0_5(N138, keyinput5, keyinput_Wire_0[5]);
not NOT1_12 (N139, N69);
  not NOT1_13 (keyinput_Wire_0[6], N76);
  xnor keyGate_0_6(KeyNOTWire_0[3], keyinput6, keyinput_Wire_0[6]);
  not KeyNOTGate_0_3(N142, KeyNOTWire_0[3]);
not NOT1_14 (N143, N82);
  not NOT1_15 (keyinput_Wire_0[7], N89);
  xor keyGate_0_7(KeyNOTWire_0[4], keyinput7, keyinput_Wire_0[7]);
  not KeyNOTGate_0_4(N146, KeyNOTWire_0[4]);
not NOT1_16 (N147, N95);
  not NOT1_17 (keyinput_Wire_0[8], N102);
  xnor keyGate_0_8(KeyNOTWire_0[5], keyinput8, keyinput_Wire_0[8]);
  not KeyNOTGate_0_5(N150, KeyNOTWire_0[5]);
not NOT1_18 (N151, N108);
  nand NAND2_19 (keyinput_Wire_0[9], N118, N4);
  xnor keyGate_0_9(KeyNOTWire_0[6], keyinput9, keyinput_Wire_0[9]);
  not KeyNOTGate_0_6(N154, KeyNOTWire_0[6]);
nor NOR2_20 (N157, N8, N119);
nor NOR2_21 (N158, N14, N119);
  nand NAND2_22 (keyinput_Wire_0[10], N122, N17);
  xor keyGate_0_10(KeyNOTWire_0[7], keyinput10, keyinput_Wire_0[10]);
  not KeyNOTGate_0_7(N159, KeyNOTWire_0[7]);
  nand NAND2_23 (keyinput_Wire_0[11], N126, N30);
  xor keyGate_0_11(KeyNOTWire_0[8], keyinput11, keyinput_Wire_0[11]);
  not KeyNOTGate_0_8(N162, KeyNOTWire_0[8]);
  nand NAND2_24 (keyinput_Wire_0[12], N130, N43);
  xnor keyGate_0_12(KeyNOTWire_0[9], keyinput12, keyinput_Wire_0[12]);
  not KeyNOTGate_0_9(N165, KeyNOTWire_0[9]);
  nand NAND2_25 (keyinput_Wire_0[13], N134, N56);
  xnor keyGate_0_13(KeyNOTWire_0[10], keyinput13, keyinput_Wire_0[13]);
  not KeyNOTGate_0_10(N168, KeyNOTWire_0[10]);
  nand NAND2_26 (keyinput_Wire_0[14], N138, N69);
  xor keyGate_0_14(KeyNOTWire_0[11], keyinput14, keyinput_Wire_0[14]);
  not KeyNOTGate_0_11(N171, KeyNOTWire_0[11]);
  nand NAND2_27 (keyinput_Wire_0[15], N142, N82);
  xnor keyGate_0_15(KeyNOTWire_0[12], keyinput15, keyinput_Wire_0[15]);
  not KeyNOTGate_0_12(N174, KeyNOTWire_0[12]);
  nand NAND2_28 (keyinput_Wire_0[16], N146, N95);
  xor keyGate_0_16(N177, keyinput16, keyinput_Wire_0[16]);
  nand NAND2_29 (keyinput_Wire_0[17], N150, N108);
  xnor keyGate_0_17(N180, keyinput17, keyinput_Wire_0[17]);
nor NOR2_30 (N183, N21, N123);
nor NOR2_31 (N184, N27, N123);
nor NOR2_32 (N185, N34, N127);
nor NOR2_33 (N186, N40, N127);
nor NOR2_34 (N187, N47, N131);
nor NOR2_35 (N188, N53, N131);
nor NOR2_36 (N189, N60, N135);
nor NOR2_37 (N190, N66, N135);
nor NOR2_38 (N191, N73, N139);
nor NOR2_39 (N192, N79, N139);
nor NOR2_40 (N193, N86, N143);
nor NOR2_41 (N194, N92, N143);
nor NOR2_42 (N195, N99, N147);
nor NOR2_43 (N196, N105, N147);
nor NOR2_44 (N197, N112, N151);
nor NOR2_45 (N198, N115, N151);
  and AND9_46 (keyinput_Wire_0[18], N154, N159, N162, N165, N168, N171, N174, N177, N180);
  xor keyGate_0_18(KeyNOTWire_0[13], keyinput18, keyinput_Wire_0[18]);
  not KeyNOTGate_0_13(N199, KeyNOTWire_0[13]);
  not NOT1_47 (keyinput_Wire_0[19], N199);
  xor keyGate_0_19(N203, keyinput19, keyinput_Wire_0[19]);
not NOT1_48 (N213, N199);
not NOT1_49 (N223, N199);
  xor XOR2_50 (keyinput_Wire_0[20], N203, N154);
  xnor keyGate_0_20(N224, keyinput20, keyinput_Wire_0[20]);
  xor XOR2_51 (keyinput_Wire_0[21], N203, N159);
  xnor keyGate_0_21(KeyNOTWire_0[14], keyinput21, keyinput_Wire_0[21]);
  not KeyNOTGate_0_14(N227, KeyNOTWire_0[14]);
  xor XOR2_52 (keyinput_Wire_0[22], N203, N162);
  xor keyGate_0_22(N230, keyinput22, keyinput_Wire_0[22]);
  xor XOR2_53 (keyinput_Wire_0[23], N203, N165);
  xnor keyGate_0_23(KeyNOTWire_0[15], keyinput23, keyinput_Wire_0[23]);
  not KeyNOTGate_0_15(N233, KeyNOTWire_0[15]);
  xor XOR2_54 (keyinput_Wire_0[24], N203, N168);
  xnor keyGate_0_24(N236, keyinput24, keyinput_Wire_0[24]);
  xor XOR2_55 (keyinput_Wire_0[25], N203, N171);
  xor keyGate_0_25(N239, keyinput25, keyinput_Wire_0[25]);
nand NAND2_56 (N242, N1, N213);
  xor XOR2_57 (keyinput_Wire_0[26], N203, N174);
  xor keyGate_0_26(N243, keyinput26, keyinput_Wire_0[26]);
nand NAND2_58 (N246, N213, N11);
xor XOR2_59 (N247, N203, N177);
nand NAND2_60 (N250, N213, N24);
  xor XOR2_61 (keyinput_Wire_0[27], N203, N180);
  xnor keyGate_0_27(N251, keyinput27, keyinput_Wire_0[27]);
nand NAND2_62 (N254, N213, N37);
nand NAND2_63 (N255, N213, N50);
nand NAND2_64 (N256, N213, N63);
nand NAND2_65 (N257, N213, N76);
nand NAND2_66 (N258, N213, N89);
nand NAND2_67 (N259, N213, N102);
nand NAND2_68 (N260, N224, N157);
nand NAND2_69 (N263, N224, N158);
nand NAND2_70 (N264, N227, N183);
nand NAND2_71 (N267, N230, N185);
nand NAND2_72 (N270, N233, N187);
nand NAND2_73 (N273, N236, N189);
nand NAND2_74 (N276, N239, N191);
nand NAND2_75 (N279, N243, N193);
nand NAND2_76 (N282, N247, N195);
nand NAND2_77 (N285, N251, N197);
nand NAND2_78 (N288, N227, N184);
nand NAND2_79 (N289, N230, N186);
nand NAND2_80 (N290, N233, N188);
nand NAND2_81 (N291, N236, N190);
nand NAND2_82 (N292, N239, N192);
nand NAND2_83 (N293, N243, N194);
nand NAND2_84 (N294, N247, N196);
nand NAND2_85 (N295, N251, N198);
  and AND9_86 (keyinput_Wire_0[28], N260, N264, N267, N270, N273, N276, N279, N282, N285);
  xor keyGate_0_28(KeyNOTWire_0[16], keyinput28, keyinput_Wire_0[28]);
  not KeyNOTGate_0_16(N296, KeyNOTWire_0[16]);
not NOT1_87 (N300, N263);
not NOT1_88 (N301, N288);
not NOT1_89 (N302, N289);
not NOT1_90 (N303, N290);
not NOT1_91 (N304, N291);
not NOT1_92 (N305, N292);
not NOT1_93 (N306, N293);
not NOT1_94 (N307, N294);
not NOT1_95 (N308, N295);
  not NOT1_96 (keyinput_Wire_0[29], N296);
  xnor keyGate_0_29(KeyNOTWire_0[17], keyinput29, keyinput_Wire_0[29]);
  not KeyNOTGate_0_17(N309, KeyNOTWire_0[17]);
not NOT1_97 (N319, N296);
not NOT1_98 (N329, N296);
xor XOR2_99 (N330, N309, N260);
xor XOR2_100 (N331, N309, N264);
xor XOR2_101 (N332, N309, N267);
xor XOR2_102 (N333, N309, N270);
nand NAND2_103 (N334, N8, N319);
xor XOR2_104 (N335, N309, N273);
nand NAND2_105 (N336, N319, N21);
xor XOR2_106 (N337, N309, N276);
nand NAND2_107 (N338, N319, N34);
xor XOR2_108 (N339, N309, N279);
nand NAND2_109 (N340, N319, N47);
xor XOR2_110 (N341, N309, N282);
nand NAND2_111 (N342, N319, N60);
xor XOR2_112 (N343, N309, N285);
nand NAND2_113 (N344, N319, N73);
nand NAND2_114 (N345, N319, N86);
nand NAND2_115 (N346, N319, N99);
nand NAND2_116 (N347, N319, N112);
nand NAND2_117 (N348, N330, N300);
nand NAND2_118 (N349, N331, N301);
nand NAND2_119 (N350, N332, N302);
nand NAND2_120 (N351, N333, N303);
nand NAND2_121 (N352, N335, N304);
nand NAND2_122 (N353, N337, N305);
nand NAND2_123 (N354, N339, N306);
nand NAND2_124 (N355, N341, N307);
nand NAND2_125 (N356, N343, N308);
  and AND9_126 (keyinput_Wire_0[30], N348, N349, N350, N351, N352, N353, N354, N355, N356);
  xnor keyGate_0_30(KeyNOTWire_0[18], keyinput30, keyinput_Wire_0[30]);
  not KeyNOTGate_0_18(N357, KeyNOTWire_0[18]);
  not NOT1_127 (keyinput_Wire_0[31], N357);
  xnor keyGate_0_31(N360, keyinput31, keyinput_Wire_0[31]);
not NOT1_128 (KeyWire_0_1, N357);
  xor flip_it (N370, KeyWire_0_1, KeyWire_0_2 );
  nand NAND2_129 (keyinput_Wire_0[32], N14, N360);
  xor keyGate_0_32(KeyNOTWire_0[19], keyinput32, keyinput_Wire_0[32]);
  not KeyNOTGate_0_19(N371, KeyNOTWire_0[19]);
  nand NAND2_130 (keyinput_Wire_0[33], N360, N27);
  xnor keyGate_0_33(N372, keyinput33, keyinput_Wire_0[33]);
  nand NAND2_131 (keyinput_Wire_0[34], N360, N40);
  xor keyGate_0_34(KeyNOTWire_0[20], keyinput34, keyinput_Wire_0[34]);
  not KeyNOTGate_0_20(N373, KeyNOTWire_0[20]);
  nand NAND2_132 (keyinput_Wire_0[35], N360, N53);
  xor keyGate_0_35(N374, keyinput35, keyinput_Wire_0[35]);
  nand NAND2_133 (keyinput_Wire_0[36], N360, N66);
  xnor keyGate_0_36(KeyNOTWire_0[21], keyinput36, keyinput_Wire_0[36]);
  not KeyNOTGate_0_21(N375, KeyNOTWire_0[21]);
  nand NAND2_134 (keyinput_Wire_0[37], N360, N79);
  xnor keyGate_0_37(N376, keyinput37, keyinput_Wire_0[37]);
  nand NAND2_135 (keyinput_Wire_0[38], N360, N92);
  xor keyGate_0_38(N377, keyinput38, keyinput_Wire_0[38]);
  nand NAND2_136 (keyinput_Wire_0[39], N360, N105);
  xor keyGate_0_39(KeyNOTWire_0[22], keyinput39, keyinput_Wire_0[39]);
  not KeyNOTGate_0_22(N378, KeyNOTWire_0[22]);
  nand NAND2_137 (keyinput_Wire_0[40], N360, N115);
  xnor keyGate_0_40(N379, keyinput40, keyinput_Wire_0[40]);
  nand NAND4_138 (keyinput_Wire_0[41], N4, N242, N334, N371);
  xor keyGate_0_41(KeyNOTWire_0[23], keyinput41, keyinput_Wire_0[41]);
  not KeyNOTGate_0_23(N380, KeyNOTWire_0[23]);
  nand NAND4_139 (keyinput_Wire_0[42], N246, N336, N372, N17);
  xor keyGate_0_42(N381, keyinput42, keyinput_Wire_0[42]);
  nand NAND4_140 (keyinput_Wire_0[43], N250, N338, N373, N30);
  xnor keyGate_0_43(N386, keyinput43, keyinput_Wire_0[43]);
  nand NAND4_141 (keyinput_Wire_0[44], N254, N340, N374, N43);
  xnor keyGate_0_44(KeyNOTWire_0[24], keyinput44, keyinput_Wire_0[44]);
  not KeyNOTGate_0_24(N393, KeyNOTWire_0[24]);
  nand NAND4_142 (keyinput_Wire_0[45], N255, N342, N375, N56);
  xnor keyGate_0_45(N399, keyinput45, keyinput_Wire_0[45]);
  nand NAND4_143 (keyinput_Wire_0[46], N256, N344, N376, N69);
  xnor keyGate_0_46(N404, keyinput46, keyinput_Wire_0[46]);
  nand NAND4_144 (keyinput_Wire_0[47], N257, N345, N377, N82);
  xnor keyGate_0_47(N407, keyinput47, keyinput_Wire_0[47]);
  nand NAND4_145 (keyinput_Wire_0[48], N258, N346, N378, N95);
  xnor keyGate_0_48(KeyNOTWire_0[25], keyinput48, keyinput_Wire_0[48]);
  not KeyNOTGate_0_25(N411, KeyNOTWire_0[25]);
  nand NAND4_146 (keyinput_Wire_0[49], N259, N347, N379, N108);
  xor keyGate_0_49(KeyNOTWire_0[26], keyinput49, keyinput_Wire_0[49]);
  not KeyNOTGate_0_26(N414, KeyNOTWire_0[26]);
  not NOT1_147 (keyinput_Wire_0[50], N380);
  xnor keyGate_0_50(KeyNOTWire_0[27], keyinput50, keyinput_Wire_0[50]);
  not KeyNOTGate_0_27(N415, KeyNOTWire_0[27]);
  and AND8_148 (keyinput_Wire_0[51], N381, N386, N393, N399, N404, N407, N411, N414);
  xnor keyGate_0_51(KeyNOTWire_0[28], keyinput51, keyinput_Wire_0[51]);
  not KeyNOTGate_0_28(N416, KeyNOTWire_0[28]);
  not NOT1_149 (keyinput_Wire_0[52], N393);
  xnor keyGate_0_52(KeyNOTWire_0[29], keyinput52, keyinput_Wire_0[52]);
  not KeyNOTGate_0_29(N417, KeyNOTWire_0[29]);
  not NOT1_150 (keyinput_Wire_0[53], N404);
  xnor keyGate_0_53(KeyNOTWire_0[30], keyinput53, keyinput_Wire_0[53]);
  not KeyNOTGate_0_30(N418, KeyNOTWire_0[30]);
  not NOT1_151 (keyinput_Wire_0[54], N407);
  xnor keyGate_0_54(KeyNOTWire_0[31], keyinput54, keyinput_Wire_0[54]);
  not KeyNOTGate_0_31(N419, KeyNOTWire_0[31]);
  not NOT1_152 (keyinput_Wire_0[55], N411);
  xnor keyGate_0_55(N420, keyinput55, keyinput_Wire_0[55]);
  nor NOR2_153 (keyinput_Wire_0[56], N415, N416);
  xnor keyGate_0_56(N421, keyinput56, keyinput_Wire_0[56]);
  nand NAND2_154 (keyinput_Wire_0[57], N386, N417);
  xor keyGate_0_57(KeyNOTWire_0[32], keyinput57, keyinput_Wire_0[57]);
  not KeyNOTGate_0_32(N422, KeyNOTWire_0[32]);
  nand NAND4_155 (keyinput_Wire_0[58], N386, N393, N418, N399);
  xor keyGate_0_58(KeyNOTWire_0[33], keyinput58, keyinput_Wire_0[58]);
  not KeyNOTGate_0_33(N425, KeyNOTWire_0[33]);
  nand NAND3_156 (keyinput_Wire_0[59], N399, N393, N419);
  xor keyGate_0_59(KeyNOTWire_0[34], keyinput59, keyinput_Wire_0[59]);
  not KeyNOTGate_0_34(N428, KeyNOTWire_0[34]);
  nand NAND4_157 (keyinput_Wire_0[60], N386, N393, N407, N420);
  xnor keyGate_0_60(KeyNOTWire_0[35], keyinput60, keyinput_Wire_0[60]);
  not KeyNOTGate_0_35(N429, KeyNOTWire_0[35]);
  nand NAND4_158 (keyinput_Wire_0[61], N381, N386, N422, N399);
  xor keyGate_0_61(KeyNOTWire_0[36], keyinput61, keyinput_Wire_0[61]);
  not KeyNOTGate_0_36(N430, KeyNOTWire_0[36]);
  nand NAND4_159 (keyinput_Wire_0[62], N381, N386, N425, N428);
  xnor keyGate_0_62(N431, keyinput62, keyinput_Wire_0[62]);
  nand NAND4_160 (keyinput_Wire_0[63], N381, N422, N425, N429);
  xnor keyGate_0_63(KeyNOTWire_0[37], keyinput63, keyinput_Wire_0[63]);
  not KeyNOTGate_0_37(N432, KeyNOTWire_0[37]);

AntiSAT some_name( KeyWire_0_2, N14, N115, N50, N105, N108, N76, N27, N47, N56, N53, N112, N63, N43, N95, N4, N34, N79, N66, N73, N40, N8, N21, N11, N102, N92, N24, N30, N69, N82, N86, N17, N37, N60, N89, N1, N99, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135,
       keyinput136, keyinput137, keyinput138, keyinput139, keyinput140,
       keyinput141, keyinput142, keyinput143, keyinput144, keyinput145,
       keyinput146, keyinput147, keyinput148, keyinput149, keyinput150,
       keyinput151, keyinput152, keyinput153, keyinput154, keyinput155,
       keyinput156, keyinput157, keyinput158, keyinput159, keyinput160,
       keyinput161, keyinput162, keyinput163, keyinput164, keyinput165,
       keyinput166, keyinput167, keyinput168, keyinput169, keyinput170,
       keyinput171);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N14, N115, N50, N105, N108, N76, N27, N47, N56, N53, N112, N63, N43, N95, N4, N34, N79, N66, N73, N40, N8, N21, N11, N102, N92, N24, N30, N69, N82, N86, N17, N37, N60, N89, N1, N99, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135 ,
        keyinput136, keyinput137, keyinput138, keyinput139, keyinput140,
        keyinput141, keyinput142, keyinput143, keyinput144, keyinput145,
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150,
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155,
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160,
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165,
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170,
        keyinput171);

  input keyinput136, keyinput137, keyinput138, keyinput139, keyinput140;
  input keyinput141, keyinput142, keyinput143, keyinput144, keyinput145;
  input keyinput146, keyinput147, keyinput148, keyinput149, keyinput150;
  input keyinput151, keyinput152, keyinput153, keyinput154, keyinput155;
  input keyinput156, keyinput157, keyinput158, keyinput159, keyinput160;
  input keyinput161, keyinput162, keyinput163, keyinput164, keyinput165;
  input keyinput166, keyinput167, keyinput168, keyinput169, keyinput170;
  input keyinput171;

  wire [0:35] keyNTin_Wire_1;
  wire [0:19] KeyNOTWire_1;

  input N14, N115, N50, N105, N108, N76, N27, N47, N56, N53, N112, N63, N43, N95, N4, N34, N79, N66, N73, N40, N8, N21, N11, N102, N92, N24, N30, N69, N82, N86, N17, N37, N60, N89, N1, N99;
  input keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73 ;

  xnor KeyGate0 (newWire_0, N14, keyinput64);
  xnor KeyGate1 (newWire_1, N115, keyinput65);
  xnor KeyGate2 (newWire_2, N50, keyinput66);
  xor  KeyGate3 (newWire_3, N105, keyinput67);
  xnor KeyGate4 (keyNTin_Wire_1[0], N108, keyinput68);
  xor keyNTinGate_1_0(newWire_4, keyinput136, keyNTin_Wire_1[0]);
  xnor KeyGate5 (keyNTin_Wire_1[1], N76, keyinput69);
  xnor keyNTinGate_1_1(newWire_5, keyinput137, keyNTin_Wire_1[1]);
  xor  KeyGate6 (newWire_6, N27, keyinput70);
  xor  KeyGate7 (keyNTin_Wire_1[2], N47, keyinput71);
  xor keyNTinGate_1_2(KeyNOTWire_1[0], keyinput138, keyNTin_Wire_1[2]);
  not KeyNOTGate_1_0(newWire_7, KeyNOTWire_1[0]);
  xor  KeyGate8 (keyNTin_Wire_1[3], N56, keyinput72);
  xor keyNTinGate_1_3(newWire_8, keyinput139, keyNTin_Wire_1[3]);
  xnor KeyGate9 (keyNTin_Wire_1[4], N53, keyinput73);
  xor keyNTinGate_1_4(KeyNOTWire_1[1], keyinput140, keyNTin_Wire_1[4]);
  not KeyNOTGate_1_1(newWire_9, KeyNOTWire_1[1]);
  xor  KeyGate10 (newWire_10, N112, keyinput74);
  xor  KeyGate11 (newWire_11, N63, keyinput75);
  xor  KeyGate12 (keyNTin_Wire_1[5], N43, keyinput76);
  xnor keyNTinGate_1_5(KeyNOTWire_1[2], keyinput141, keyNTin_Wire_1[5]);
  not KeyNOTGate_1_2(newWire_12, KeyNOTWire_1[2]);
  xnor KeyGate13 (newWire_13, N95, keyinput77);
  xnor KeyGate14 (newWire_14, N4, keyinput78);
  xnor KeyGate15 (keyNTin_Wire_1[6], N34, keyinput79);
  xor keyNTinGate_1_6(KeyNOTWire_1[3], keyinput142, keyNTin_Wire_1[6]);
  not KeyNOTGate_1_3(newWire_15, KeyNOTWire_1[3]);
  xor  KeyGate16 (newWire_16, N79, keyinput80);
  xor  KeyGate17 (newWire_17, N66, keyinput81);
  xnor KeyGate18 (newWire_18, N73, keyinput82);
  xnor KeyGate19 (keyNTin_Wire_1[7], N40, keyinput83);
  xnor keyNTinGate_1_7(KeyNOTWire_1[4], keyinput143, keyNTin_Wire_1[7]);
  not KeyNOTGate_1_4(newWire_19, KeyNOTWire_1[4]);
  xor  KeyGate20 (newWire_20, N8, keyinput84);
  xor  KeyGate21 (keyNTin_Wire_1[8], N21, keyinput85);
  xor keyNTinGate_1_8(newWire_21, keyinput144, keyNTin_Wire_1[8]);
  xnor KeyGate22 (keyNTin_Wire_1[9], N11, keyinput86);
  xor keyNTinGate_1_9(newWire_22, keyinput145, keyNTin_Wire_1[9]);
  xor  KeyGate23 (newWire_23, N102, keyinput87);
  xnor KeyGate24 (keyNTin_Wire_1[10], N92, keyinput88);
  xor keyNTinGate_1_10(newWire_24, keyinput146, keyNTin_Wire_1[10]);
  xnor KeyGate25 (keyNTin_Wire_1[11], N24, keyinput89);
  xor keyNTinGate_1_11(KeyNOTWire_1[5], keyinput147, keyNTin_Wire_1[11]);
  not KeyNOTGate_1_5(newWire_25, KeyNOTWire_1[5]);
  xnor KeyGate26 (newWire_26, N30, keyinput90);
  xor  KeyGate27 (newWire_27, N69, keyinput91);
  xnor KeyGate28 (keyNTin_Wire_1[12], N82, keyinput92);
  xor keyNTinGate_1_12(newWire_28, keyinput148, keyNTin_Wire_1[12]);
  xor  KeyGate29 (newWire_29, N86, keyinput93);
  xor  KeyGate30 (newWire_30, N17, keyinput94);
  xor  KeyGate31 (keyNTin_Wire_1[13], N37, keyinput95);
  xnor keyNTinGate_1_13(KeyNOTWire_1[6], keyinput149, keyNTin_Wire_1[13]);
  not KeyNOTGate_1_6(newWire_31, KeyNOTWire_1[6]);
  xnor KeyGate32 (keyNTin_Wire_1[14], N60, keyinput96);
  xnor keyNTinGate_1_14(KeyNOTWire_1[7], keyinput150, keyNTin_Wire_1[14]);
  not KeyNOTGate_1_7(newWire_32, KeyNOTWire_1[7]);
  xor  KeyGate33 (keyNTin_Wire_1[15], N89, keyinput97);
  xnor keyNTinGate_1_15(KeyNOTWire_1[8], keyinput151, keyNTin_Wire_1[15]);
  not KeyNOTGate_1_8(newWire_33, KeyNOTWire_1[8]);
  xnor KeyGate34 (newWire_34, N1, keyinput98);
  xnor KeyGate35 (keyNTin_Wire_1[16], N99, keyinput99);
  xnor keyNTinGate_1_16(newWire_35, keyinput152, keyNTin_Wire_1[16]);
  xnor KeyGate36 (newWire_36, N14, keyinput100);
  xor  KeyGate37 (newWire_37, N115, keyinput101);
  xor  KeyGate38 (newWire_38, N50, keyinput102);
  xor  KeyGate39 (keyNTin_Wire_1[17], N105, keyinput103);
  xnor keyNTinGate_1_17(newWire_39, keyinput153, keyNTin_Wire_1[17]);
  xor  KeyGate40 (newWire_40, N108, keyinput104);
  xor  KeyGate41 (newWire_41, N76, keyinput105);
  xnor KeyGate42 (newWire_42, N27, keyinput106);
  xnor KeyGate43 (keyNTin_Wire_1[18], N47, keyinput107);
  xor keyNTinGate_1_18(KeyNOTWire_1[9], keyinput154, keyNTin_Wire_1[18]);
  not KeyNOTGate_1_9(newWire_43, KeyNOTWire_1[9]);
  xor  KeyGate44 (keyNTin_Wire_1[19], N56, keyinput108);
  xor keyNTinGate_1_19(KeyNOTWire_1[10], keyinput155, keyNTin_Wire_1[19]);
  not KeyNOTGate_1_10(newWire_44, KeyNOTWire_1[10]);
  xnor KeyGate45 (newWire_45, N53, keyinput109);
  xor  KeyGate46 (keyNTin_Wire_1[20], N112, keyinput110);
  xnor keyNTinGate_1_20(newWire_46, keyinput156, keyNTin_Wire_1[20]);
  xor  KeyGate47 (newWire_47, N63, keyinput111);
  xor  KeyGate48 (keyNTin_Wire_1[21], N43, keyinput112);
  xor keyNTinGate_1_21(KeyNOTWire_1[11], keyinput157, keyNTin_Wire_1[21]);
  not KeyNOTGate_1_11(newWire_48, KeyNOTWire_1[11]);
  xnor KeyGate49 (newWire_49, N95, keyinput113);
  xor  KeyGate50 (newWire_50, N4, keyinput114);
  xnor KeyGate51 (keyNTin_Wire_1[22], N34, keyinput115);
  xor keyNTinGate_1_22(KeyNOTWire_1[12], keyinput158, keyNTin_Wire_1[22]);
  not KeyNOTGate_1_12(newWire_51, KeyNOTWire_1[12]);
  xnor KeyGate52 (keyNTin_Wire_1[23], N79, keyinput116);
  xnor keyNTinGate_1_23(KeyNOTWire_1[13], keyinput159, keyNTin_Wire_1[23]);
  not KeyNOTGate_1_13(newWire_52, KeyNOTWire_1[13]);
  xnor KeyGate53 (keyNTin_Wire_1[24], N66, keyinput117);
  xor keyNTinGate_1_24(newWire_53, keyinput160, keyNTin_Wire_1[24]);
  xor  KeyGate54 (newWire_54, N73, keyinput118);
  xor  KeyGate55 (keyNTin_Wire_1[25], N40, keyinput119);
  xor keyNTinGate_1_25(newWire_55, keyinput161, keyNTin_Wire_1[25]);
  xnor KeyGate56 (newWire_56, N8, keyinput120);
  xor  KeyGate57 (keyNTin_Wire_1[26], N21, keyinput121);
  xnor keyNTinGate_1_26(KeyNOTWire_1[14], keyinput162, keyNTin_Wire_1[26]);
  not KeyNOTGate_1_14(newWire_57, KeyNOTWire_1[14]);
  xor  KeyGate58 (newWire_58, N11, keyinput122);
  xor  KeyGate59 (newWire_59, N102, keyinput123);
  xor  KeyGate60 (newWire_60, N92, keyinput124);
  xnor KeyGate61 (keyNTin_Wire_1[27], N24, keyinput125);
  xor keyNTinGate_1_27(KeyNOTWire_1[15], keyinput163, keyNTin_Wire_1[27]);
  not KeyNOTGate_1_15(newWire_61, KeyNOTWire_1[15]);
  xnor KeyGate62 (keyNTin_Wire_1[28], N30, keyinput126);
  xor keyNTinGate_1_28(newWire_62, keyinput164, keyNTin_Wire_1[28]);
  xor  KeyGate63 (newWire_63, N69, keyinput127);
  xnor KeyGate64 (keyNTin_Wire_1[29], N82, keyinput128);
  xnor keyNTinGate_1_29(newWire_64, keyinput165, keyNTin_Wire_1[29]);
  xor  KeyGate65 (keyNTin_Wire_1[30], N86, keyinput129);
  xor keyNTinGate_1_30(KeyNOTWire_1[16], keyinput166, keyNTin_Wire_1[30]);
  not KeyNOTGate_1_16(newWire_65, KeyNOTWire_1[16]);
  xnor KeyGate66 (keyNTin_Wire_1[31], N17, keyinput130);
  xnor keyNTinGate_1_31(KeyNOTWire_1[17], keyinput167, keyNTin_Wire_1[31]);
  not KeyNOTGate_1_17(newWire_66, KeyNOTWire_1[17]);
  xnor KeyGate67 (newWire_67, N37, keyinput131);
  xnor KeyGate68 (keyNTin_Wire_1[32], N60, keyinput132);
  xnor keyNTinGate_1_32(KeyNOTWire_1[18], keyinput168, keyNTin_Wire_1[32]);
  not KeyNOTGate_1_18(newWire_68, KeyNOTWire_1[18]);
  xor  KeyGate69 (newWire_69, N89, keyinput133);
  xor  KeyGate70 (newWire_70, N1, keyinput134);
  xnor KeyGate71 (keyNTin_Wire_1[33], N99, keyinput135);
  xor keyNTinGate_1_33(newWire_71, keyinput169, keyNTin_Wire_1[33]);
  and some_function (keyNTin_Wire_1[34], newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35 );
  xor keyNTinGate_1_34(KeyNOTWire_1[19], keyinput170, keyNTin_Wire_1[34]);
  not KeyNOTGate_1_19(newWire_72, KeyNOTWire_1[19]);
  nand compl_function (keyNTin_Wire_1[35], newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71);
  xnor keyNTinGate_1_35(newWire_73, keyinput171, keyNTin_Wire_1[35]);
  and finalAND (KeyWire_0_2, newWire_72, newWire_73);

endmodule /* AntiSAT */
