`timescale 1ns / 1ps
// Verilog
// c880
// Ninputs 60
// Noutputs 26
// NtotalGates 383
// NAND4 13
// AND3 12
// NAND2 60
// NAND3 14
// AND2 105
// OR2 29
// NOT1 63
// NOR2 61
// BUFF1 26

module top (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
                  N865,N866,N874,N878,N879,N880,
        keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4,
        keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9,
        keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14,
        keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19,
        keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24,
        keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29,
        keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34,
        keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39,
        keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44,
        keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49,
        keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54,
        keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59,
        keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64,
        keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69,
        keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74,
        keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79,
        keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84,
        keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89,
        keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94,
        keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99,
        keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104,
        keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109,
        keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114,
        keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119,
        keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124,
        keyIn_0_125, keyIn_0_126, keyIn_0_127);

  input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4;
  input keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9;
  input keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14;
  input keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19;
  input keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24;
  input keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29;
  input keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34;
  input keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39;
  input keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44;
  input keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49;
  input keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54;
  input keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59;
  input keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64;
  input keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69;
  input keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74;
  input keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79;
  input keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84;
  input keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89;
  input keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94;
  input keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99;
  input keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104;
  input keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109;
  input keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114;
  input keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119;
  input keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124;
  input keyIn_0_125, keyIn_0_126, keyIn_0_127;

  wire [0:127] KeyWire_0;
  wire [0:54] KeyNOTWire_0;

input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;

output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;

wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877;

nand NAND4_1 (N269, N1, N8, N13, N17);
nand NAND4_2 (N270, N1, N26, N13, N17);
and AND3_3 (N273, N29, N36, N42);
  and AND3_4 (KeyWire_0[0], N1, N26, N51);
  xor KeyGate_0_0(N276, keyIn_0_0, KeyWire_0[0]);
  nand NAND4_5 (KeyWire_0[1], N1, N8, N51, N17);
  xnor KeyGate_0_1(N279, keyIn_0_1, KeyWire_0[1]);
nand NAND4_6 (N280, N1, N8, N13, N55);
nand NAND4_7 (N284, N59, N42, N68, N72);
nand NAND2_8 (N285, N29, N68);
nand NAND3_9 (N286, N59, N68, N74);
  and AND3_10 (KeyWire_0[2], N29, N75, N80);
  xor KeyGate_0_2(KeyNOTWire_0[0], keyIn_0_2, KeyWire_0[2]);
  not KeyNOTGate_0_0(N287, KeyNOTWire_0[0]);
and AND3_11 (N290, N29, N75, N42);
and AND3_12 (N291, N29, N36, N80);
and AND3_13 (N292, N29, N36, N42);
and AND3_14 (N293, N59, N75, N80);
  and AND3_15 (KeyWire_0[3], N59, N75, N42);
  xnor KeyGate_0_3(N294, keyIn_0_3, KeyWire_0[3]);
and AND3_16 (N295, N59, N36, N80);
and AND3_17 (N296, N59, N36, N42);
and AND2_18 (N297, N85, N86);
or OR2_19 (N298, N87, N88);
nand NAND2_20 (N301, N91, N96);
or OR2_21 (N302, N91, N96);
nand NAND2_22 (N303, N101, N106);
or OR2_23 (N304, N101, N106);
nand NAND2_24 (N305, N111, N116);
or OR2_25 (N306, N111, N116);
nand NAND2_26 (N307, N121, N126);
or OR2_27 (N308, N121, N126);
and AND2_28 (N309, N8, N138);
  not NOT1_29 (KeyWire_0[4], N268);
  xnor KeyGate_0_4(N310, keyIn_0_4, KeyWire_0[4]);
and AND2_30 (N316, N51, N138);
and AND2_31 (N317, N17, N138);
and AND2_32 (N318, N152, N138);
  nand NAND2_33 (KeyWire_0[5], N59, N156);
  xnor KeyGate_0_5(N319, keyIn_0_5, KeyWire_0[5]);
  nor NOR2_34 (KeyWire_0[6], N17, N42);
  xor KeyGate_0_6(N322, keyIn_0_6, KeyWire_0[6]);
  and AND2_35 (KeyWire_0[7], N17, N42);
  xor KeyGate_0_7(N323, keyIn_0_7, KeyWire_0[7]);
nand NAND2_36 (N324, N159, N165);
or OR2_37 (N325, N159, N165);
nand NAND2_38 (N326, N171, N177);
or OR2_39 (N327, N171, N177);
nand NAND2_40 (N328, N183, N189);
or OR2_41 (N329, N183, N189);
nand NAND2_42 (N330, N195, N201);
or OR2_43 (N331, N195, N201);
and AND2_44 (N332, N210, N91);
and AND2_45 (N333, N210, N96);
and AND2_46 (N334, N210, N101);
and AND2_47 (N335, N210, N106);
and AND2_48 (N336, N210, N111);
and AND2_49 (N337, N255, N259);
and AND2_50 (N338, N210, N116);
and AND2_51 (N339, N255, N260);
and AND2_52 (N340, N210, N121);
and AND2_53 (N341, N255, N267);
not NOT1_54 (N342, N269);
not NOT1_55 (N343, N273);
or OR2_56 (N344, N270, N273);
  not NOT1_57 (KeyWire_0[8], N276);
  xor KeyGate_0_8(N345, keyIn_0_8, KeyWire_0[8]);
not NOT1_58 (N346, N276);
  not NOT1_59 (KeyWire_0[9], N279);
  xor KeyGate_0_9(KeyNOTWire_0[1], keyIn_0_9, KeyWire_0[9]);
  not KeyNOTGate_0_1(N347, KeyNOTWire_0[1]);
nor NOR2_60 (N348, N280, N284);
or OR2_61 (N349, N280, N285);
  or OR2_62 (KeyWire_0[10], N280, N286);
  xnor KeyGate_0_10(KeyNOTWire_0[2], keyIn_0_10, KeyWire_0[10]);
  not KeyNOTGate_0_2(N350, KeyNOTWire_0[2]);
not NOT1_63 (N351, N293);
  not NOT1_64 (KeyWire_0[11], N294);
  xnor KeyGate_0_11(N352, keyIn_0_11, KeyWire_0[11]);
not NOT1_65 (N353, N295);
not NOT1_66 (N354, N296);
nand NAND2_67 (N355, N89, N298);
and AND2_68 (N356, N90, N298);
nand NAND2_69 (N357, N301, N302);
nand NAND2_70 (N360, N303, N304);
nand NAND2_71 (N363, N305, N306);
nand NAND2_72 (N366, N307, N308);
  not NOT1_73 (KeyWire_0[12], N310);
  xnor KeyGate_0_12(N369, keyIn_0_12, KeyWire_0[12]);
  nor NOR2_74 (KeyWire_0[13], N322, N323);
  xor KeyGate_0_13(KeyNOTWire_0[3], keyIn_0_13, KeyWire_0[13]);
  not KeyNOTGate_0_3(N375, KeyNOTWire_0[3]);
nand NAND2_75 (N376, N324, N325);
nand NAND2_76 (N379, N326, N327);
nand NAND2_77 (N382, N328, N329);
nand NAND2_78 (N385, N330, N331);
buf BUFF1_79 (N388, N290);
buf BUFF1_80 (N389, N291);
buf BUFF1_81 (N390, N292);
buf BUFF1_82 (N391, N297);
or OR2_83 (N392, N270, N343);
  not NOT1_84 (KeyWire_0[14], N345);
  xor KeyGate_0_14(N393, keyIn_0_14, KeyWire_0[14]);
not NOT1_85 (N399, N346);
and AND2_86 (N400, N348, N73);
not NOT1_87 (N401, N349);
not NOT1_88 (N402, N350);
not NOT1_89 (N403, N355);
not NOT1_90 (N404, N357);
  not NOT1_91 (KeyWire_0[15], N360);
  xnor KeyGate_0_15(N405, keyIn_0_15, KeyWire_0[15]);
and AND2_92 (N406, N357, N360);
not NOT1_93 (N407, N363);
not NOT1_94 (N408, N366);
and AND2_95 (N409, N363, N366);
  nand NAND2_96 (KeyWire_0[16], N347, N352);
  xnor KeyGate_0_16(KeyNOTWire_0[4], keyIn_0_16, KeyWire_0[16]);
  not KeyNOTGate_0_4(N410, KeyNOTWire_0[4]);
not NOT1_97 (N411, N376);
not NOT1_98 (N412, N379);
and AND2_99 (N413, N376, N379);
not NOT1_100 (N414, N382);
not NOT1_101 (N415, N385);
and AND2_102 (N416, N382, N385);
and AND2_103 (N417, N210, N369);
buf BUFF1_104 (N418, N342);
buf BUFF1_105 (N419, N344);
buf BUFF1_106 (N420, N351);
buf BUFF1_107 (N421, N353);
buf BUFF1_108 (N422, N354);
buf BUFF1_109 (N423, N356);
not NOT1_110 (N424, N400);
and AND2_111 (N425, N404, N405);
and AND2_112 (N426, N407, N408);
  and AND3_113 (KeyWire_0[17], N319, N393, N55);
  xor KeyGate_0_17(KeyNOTWire_0[5], keyIn_0_17, KeyWire_0[17]);
  not KeyNOTGate_0_5(N427, KeyNOTWire_0[5]);
  and AND3_114 (KeyWire_0[18], N393, N17, N287);
  xor KeyGate_0_18(N432, keyIn_0_18, KeyWire_0[18]);
  nand NAND3_115 (KeyWire_0[19], N393, N287, N55);
  xnor KeyGate_0_19(KeyNOTWire_0[6], keyIn_0_19, KeyWire_0[19]);
  not KeyNOTGate_0_6(N437, KeyNOTWire_0[6]);
  nand NAND4_116 (KeyWire_0[20], N375, N59, N156, N393);
  xnor KeyGate_0_20(KeyNOTWire_0[7], keyIn_0_20, KeyWire_0[20]);
  not KeyNOTGate_0_7(N442, KeyNOTWire_0[7]);
  nand NAND3_117 (KeyWire_0[21], N393, N319, N17);
  xor KeyGate_0_21(KeyNOTWire_0[8], keyIn_0_21, KeyWire_0[21]);
  not KeyNOTGate_0_8(N443, KeyNOTWire_0[8]);
and AND2_118 (N444, N411, N412);
and AND2_119 (N445, N414, N415);
buf BUFF1_120 (N446, N392);
buf BUFF1_121 (N447, N399);
buf BUFF1_122 (N448, N401);
buf BUFF1_123 (N449, N402);
buf BUFF1_124 (N450, N403);
not NOT1_125 (N451, N424);
nor NOR2_126 (N460, N406, N425);
nor NOR2_127 (N463, N409, N426);
  nand NAND2_128 (KeyWire_0[22], N442, N410);
  xor KeyGate_0_22(KeyNOTWire_0[9], keyIn_0_22, KeyWire_0[22]);
  not KeyNOTGate_0_9(N466, KeyNOTWire_0[9]);
and AND2_129 (N475, N143, N427);
and AND2_130 (N476, N310, N432);
and AND2_131 (N477, N146, N427);
and AND2_132 (N478, N310, N432);
and AND2_133 (N479, N149, N427);
and AND2_134 (N480, N310, N432);
  and AND2_135 (KeyWire_0[23], N153, N427);
  xor KeyGate_0_23(KeyNOTWire_0[10], keyIn_0_23, KeyWire_0[23]);
  not KeyNOTGate_0_10(N481, KeyNOTWire_0[10]);
  and AND2_136 (KeyWire_0[24], N310, N432);
  xnor KeyGate_0_24(N482, keyIn_0_24, KeyWire_0[24]);
  nand NAND2_137 (KeyWire_0[25], N443, N1);
  xnor KeyGate_0_25(N483, keyIn_0_25, KeyWire_0[25]);
  or OR2_138 (KeyWire_0[26], N369, N437);
  xor KeyGate_0_26(N488, keyIn_0_26, KeyWire_0[26]);
  or OR2_139 (KeyWire_0[27], N369, N437);
  xnor KeyGate_0_27(N489, keyIn_0_27, KeyWire_0[27]);
  or OR2_140 (KeyWire_0[28], N369, N437);
  xor KeyGate_0_28(N490, keyIn_0_28, KeyWire_0[28]);
  or OR2_141 (KeyWire_0[29], N369, N437);
  xnor KeyGate_0_29(N491, keyIn_0_29, KeyWire_0[29]);
nor NOR2_142 (N492, N413, N444);
nor NOR2_143 (N495, N416, N445);
nand NAND2_144 (N498, N130, N460);
or OR2_145 (N499, N130, N460);
nand NAND2_146 (N500, N463, N135);
or OR2_147 (N501, N463, N135);
and AND2_148 (N502, N91, N466);
nor NOR2_149 (N503, N475, N476);
and AND2_150 (N504, N96, N466);
nor NOR2_151 (N505, N477, N478);
and AND2_152 (N506, N101, N466);
nor NOR2_153 (N507, N479, N480);
  and AND2_154 (KeyWire_0[30], N106, N466);
  xnor KeyGate_0_30(N508, keyIn_0_30, KeyWire_0[30]);
  nor NOR2_155 (KeyWire_0[31], N481, N482);
  xnor KeyGate_0_31(N509, keyIn_0_31, KeyWire_0[31]);
  and AND2_156 (KeyWire_0[32], N143, N483);
  xnor KeyGate_0_32(N510, keyIn_0_32, KeyWire_0[32]);
  and AND2_157 (KeyWire_0[33], N111, N466);
  xor KeyGate_0_33(N511, keyIn_0_33, KeyWire_0[33]);
  and AND2_158 (KeyWire_0[34], N146, N483);
  xor KeyGate_0_34(N512, keyIn_0_34, KeyWire_0[34]);
  and AND2_159 (KeyWire_0[35], N116, N466);
  xor KeyGate_0_35(N513, keyIn_0_35, KeyWire_0[35]);
  and AND2_160 (KeyWire_0[36], N149, N483);
  xor KeyGate_0_36(KeyNOTWire_0[11], keyIn_0_36, KeyWire_0[36]);
  not KeyNOTGate_0_11(N514, KeyNOTWire_0[11]);
  and AND2_161 (KeyWire_0[37], N121, N466);
  xor KeyGate_0_37(KeyNOTWire_0[12], keyIn_0_37, KeyWire_0[37]);
  not KeyNOTGate_0_12(N515, KeyNOTWire_0[12]);
  and AND2_162 (KeyWire_0[38], N153, N483);
  xnor KeyGate_0_38(KeyNOTWire_0[13], keyIn_0_38, KeyWire_0[38]);
  not KeyNOTGate_0_13(N516, KeyNOTWire_0[13]);
  and AND2_163 (KeyWire_0[39], N126, N466);
  xnor KeyGate_0_39(N517, keyIn_0_39, KeyWire_0[39]);
nand NAND2_164 (N518, N130, N492);
or OR2_165 (N519, N130, N492);
nand NAND2_166 (N520, N495, N207);
or OR2_167 (N521, N495, N207);
and AND2_168 (N522, N451, N159);
and AND2_169 (N523, N451, N165);
and AND2_170 (N524, N451, N171);
and AND2_171 (N525, N451, N177);
and AND2_172 (N526, N451, N183);
nand NAND2_173 (N527, N451, N189);
nand NAND2_174 (N528, N451, N195);
nand NAND2_175 (N529, N451, N201);
nand NAND2_176 (N530, N498, N499);
nand NAND2_177 (N533, N500, N501);
  nor NOR2_178 (KeyWire_0[40], N309, N502);
  xnor KeyGate_0_40(KeyNOTWire_0[14], keyIn_0_40, KeyWire_0[40]);
  not KeyNOTGate_0_14(N536, KeyNOTWire_0[14]);
nor NOR2_179 (N537, N316, N504);
nor NOR2_180 (N538, N317, N506);
  nor NOR2_181 (KeyWire_0[41], N318, N508);
  xnor KeyGate_0_41(N539, keyIn_0_41, KeyWire_0[41]);
  nor NOR2_182 (KeyWire_0[42], N510, N511);
  xor KeyGate_0_42(N540, keyIn_0_42, KeyWire_0[42]);
  nor NOR2_183 (KeyWire_0[43], N512, N513);
  xor KeyGate_0_43(KeyNOTWire_0[15], keyIn_0_43, KeyWire_0[43]);
  not KeyNOTGate_0_15(N541, KeyNOTWire_0[15]);
  nor NOR2_184 (KeyWire_0[44], N514, N515);
  xnor KeyGate_0_44(KeyNOTWire_0[16], keyIn_0_44, KeyWire_0[44]);
  not KeyNOTGate_0_16(N542, KeyNOTWire_0[16]);
  nor NOR2_185 (KeyWire_0[45], N516, N517);
  xor KeyGate_0_45(N543, keyIn_0_45, KeyWire_0[45]);
nand NAND2_186 (N544, N518, N519);
nand NAND2_187 (N547, N520, N521);
not NOT1_188 (N550, N530);
not NOT1_189 (N551, N533);
and AND2_190 (N552, N530, N533);
nand NAND2_191 (N553, N536, N503);
nand NAND2_192 (N557, N537, N505);
nand NAND2_193 (N561, N538, N507);
  nand NAND2_194 (KeyWire_0[46], N539, N509);
  xnor KeyGate_0_46(N565, keyIn_0_46, KeyWire_0[46]);
  nand NAND2_195 (KeyWire_0[47], N488, N540);
  xnor KeyGate_0_47(KeyNOTWire_0[17], keyIn_0_47, KeyWire_0[47]);
  not KeyNOTGate_0_17(N569, KeyNOTWire_0[17]);
  nand NAND2_196 (KeyWire_0[48], N489, N541);
  xnor KeyGate_0_48(N573, keyIn_0_48, KeyWire_0[48]);
  nand NAND2_197 (KeyWire_0[49], N490, N542);
  xor KeyGate_0_49(KeyNOTWire_0[18], keyIn_0_49, KeyWire_0[49]);
  not KeyNOTGate_0_18(N577, KeyNOTWire_0[18]);
  nand NAND2_198 (KeyWire_0[50], N491, N543);
  xnor KeyGate_0_50(N581, keyIn_0_50, KeyWire_0[50]);
not NOT1_199 (N585, N544);
not NOT1_200 (N586, N547);
and AND2_201 (N587, N544, N547);
and AND2_202 (N588, N550, N551);
and AND2_203 (N589, N585, N586);
  nand NAND2_204 (KeyWire_0[51], N553, N159);
  xor KeyGate_0_51(N590, keyIn_0_51, KeyWire_0[51]);
or OR2_205 (N593, N553, N159);
and AND2_206 (N596, N246, N553);
nand NAND2_207 (N597, N557, N165);
or OR2_208 (N600, N557, N165);
and AND2_209 (N605, N246, N557);
nand NAND2_210 (N606, N561, N171);
or OR2_211 (N609, N561, N171);
and AND2_212 (N615, N246, N561);
  nand NAND2_213 (KeyWire_0[52], N565, N177);
  xor KeyGate_0_52(KeyNOTWire_0[19], keyIn_0_52, KeyWire_0[52]);
  not KeyNOTGate_0_19(N616, KeyNOTWire_0[19]);
  or OR2_214 (KeyWire_0[53], N565, N177);
  xnor KeyGate_0_53(KeyNOTWire_0[20], keyIn_0_53, KeyWire_0[53]);
  not KeyNOTGate_0_20(N619, KeyNOTWire_0[20]);
and AND2_215 (N624, N246, N565);
  nand NAND2_216 (KeyWire_0[54], N569, N183);
  xor KeyGate_0_54(KeyNOTWire_0[21], keyIn_0_54, KeyWire_0[54]);
  not KeyNOTGate_0_21(N625, KeyNOTWire_0[21]);
  or OR2_217 (KeyWire_0[55], N569, N183);
  xor KeyGate_0_55(N628, keyIn_0_55, KeyWire_0[55]);
and AND2_218 (N631, N246, N569);
  nand NAND2_219 (KeyWire_0[56], N573, N189);
  xor KeyGate_0_56(N632, keyIn_0_56, KeyWire_0[56]);
  or OR2_220 (KeyWire_0[57], N573, N189);
  xor KeyGate_0_57(KeyNOTWire_0[22], keyIn_0_57, KeyWire_0[57]);
  not KeyNOTGate_0_22(N635, KeyNOTWire_0[22]);
and AND2_221 (N640, N246, N573);
  nand NAND2_222 (KeyWire_0[58], N577, N195);
  xor KeyGate_0_58(KeyNOTWire_0[23], keyIn_0_58, KeyWire_0[58]);
  not KeyNOTGate_0_23(N641, KeyNOTWire_0[23]);
  or OR2_223 (KeyWire_0[59], N577, N195);
  xor KeyGate_0_59(KeyNOTWire_0[24], keyIn_0_59, KeyWire_0[59]);
  not KeyNOTGate_0_24(N644, KeyNOTWire_0[24]);
and AND2_224 (N650, N246, N577);
  nand NAND2_225 (KeyWire_0[60], N581, N201);
  xnor KeyGate_0_60(N651, keyIn_0_60, KeyWire_0[60]);
  or OR2_226 (KeyWire_0[61], N581, N201);
  xnor KeyGate_0_61(N654, keyIn_0_61, KeyWire_0[61]);
and AND2_227 (N659, N246, N581);
nor NOR2_228 (N660, N552, N588);
nor NOR2_229 (N661, N587, N589);
not NOT1_230 (N662, N590);
  and AND2_231 (KeyWire_0[62], N593, N590);
  xnor KeyGate_0_62(N665, keyIn_0_62, KeyWire_0[62]);
nor NOR2_232 (N669, N596, N522);
not NOT1_233 (N670, N597);
and AND2_234 (N673, N600, N597);
nor NOR2_235 (N677, N605, N523);
not NOT1_236 (N678, N606);
and AND2_237 (N682, N609, N606);
nor NOR2_238 (N686, N615, N524);
  not NOT1_239 (KeyWire_0[63], N616);
  xor KeyGate_0_63(N687, keyIn_0_63, KeyWire_0[63]);
and AND2_240 (N692, N619, N616);
nor NOR2_241 (N696, N624, N525);
  not NOT1_242 (KeyWire_0[64], N625);
  xor KeyGate_0_64(N697, keyIn_0_64, KeyWire_0[64]);
and AND2_243 (N700, N628, N625);
nor NOR2_244 (N704, N631, N526);
  not NOT1_245 (KeyWire_0[65], N632);
  xnor KeyGate_0_65(N705, keyIn_0_65, KeyWire_0[65]);
and AND2_246 (N708, N635, N632);
nor NOR2_247 (N712, N337, N640);
  not NOT1_248 (KeyWire_0[66], N641);
  xor KeyGate_0_66(N713, keyIn_0_66, KeyWire_0[66]);
and AND2_249 (N717, N644, N641);
nor NOR2_250 (N721, N339, N650);
  not NOT1_251 (KeyWire_0[67], N651);
  xnor KeyGate_0_67(N722, keyIn_0_67, KeyWire_0[67]);
and AND2_252 (N727, N654, N651);
nor NOR2_253 (N731, N341, N659);
nand NAND2_254 (N732, N654, N261);
nand NAND3_255 (N733, N644, N654, N261);
  nand NAND4_256 (KeyWire_0[68], N635, N644, N654, N261);
  xnor KeyGate_0_68(KeyNOTWire_0[25], keyIn_0_68, KeyWire_0[68]);
  not KeyNOTGate_0_25(N734, KeyNOTWire_0[25]);
not NOT1_257 (N735, N662);
and AND2_258 (N736, N228, N665);
and AND2_259 (N737, N237, N662);
not NOT1_260 (N738, N670);
and AND2_261 (N739, N228, N673);
and AND2_262 (N740, N237, N670);
not NOT1_263 (N741, N678);
and AND2_264 (N742, N228, N682);
and AND2_265 (N743, N237, N678);
not NOT1_266 (N744, N687);
and AND2_267 (N745, N228, N692);
  and AND2_268 (KeyWire_0[69], N237, N687);
  xor KeyGate_0_69(N746, keyIn_0_69, KeyWire_0[69]);
  not NOT1_269 (KeyWire_0[70], N697);
  xnor KeyGate_0_70(KeyNOTWire_0[26], keyIn_0_70, KeyWire_0[70]);
  not KeyNOTGate_0_26(N747, KeyNOTWire_0[26]);
and AND2_270 (N748, N228, N700);
and AND2_271 (N749, N237, N697);
  not NOT1_272 (KeyWire_0[71], N705);
  xnor KeyGate_0_71(KeyNOTWire_0[27], keyIn_0_71, KeyWire_0[71]);
  not KeyNOTGate_0_27(N750, KeyNOTWire_0[27]);
and AND2_273 (N751, N228, N708);
and AND2_274 (N752, N237, N705);
not NOT1_275 (N753, N713);
and AND2_276 (N754, N228, N717);
and AND2_277 (N755, N237, N713);
not NOT1_278 (N756, N722);
nor NOR2_279 (N757, N727, N261);
and AND2_280 (N758, N727, N261);
and AND2_281 (N759, N228, N727);
and AND2_282 (N760, N237, N722);
nand NAND2_283 (N761, N644, N722);
  nand NAND2_284 (KeyWire_0[72], N635, N713);
  xnor KeyGate_0_72(N762, keyIn_0_72, KeyWire_0[72]);
  nand NAND3_285 (KeyWire_0[73], N635, N644, N722);
  xor KeyGate_0_73(KeyNOTWire_0[28], keyIn_0_73, KeyWire_0[73]);
  not KeyNOTGate_0_28(N763, KeyNOTWire_0[28]);
nand NAND2_286 (N764, N609, N687);
nand NAND2_287 (N765, N600, N678);
  nand NAND3_288 (KeyWire_0[74], N600, N609, N687);
  xor KeyGate_0_74(KeyNOTWire_0[29], keyIn_0_74, KeyWire_0[74]);
  not KeyNOTGate_0_29(N766, KeyNOTWire_0[29]);
buf BUFF1_289 (N767, N660);
buf BUFF1_290 (N768, N661);
nor NOR2_291 (N769, N736, N737);
nor NOR2_292 (N770, N739, N740);
nor NOR2_293 (N771, N742, N743);
nor NOR2_294 (N772, N745, N746);
  nand NAND4_295 (KeyWire_0[75], N750, N762, N763, N734);
  xor KeyGate_0_75(KeyNOTWire_0[30], keyIn_0_75, KeyWire_0[75]);
  not KeyNOTGate_0_30(N773, KeyNOTWire_0[30]);
nor NOR2_296 (N777, N748, N749);
nand NAND3_297 (N778, N753, N761, N733);
nor NOR2_298 (N781, N751, N752);
nand NAND2_299 (N782, N756, N732);
nor NOR2_300 (N785, N754, N755);
nor NOR2_301 (N786, N757, N758);
nor NOR2_302 (N787, N759, N760);
  nor NOR2_303 (KeyWire_0[76], N700, N773);
  xnor KeyGate_0_76(N788, keyIn_0_76, KeyWire_0[76]);
  and AND2_304 (KeyWire_0[77], N700, N773);
  xnor KeyGate_0_77(N789, keyIn_0_77, KeyWire_0[77]);
nor NOR2_305 (N790, N708, N778);
and AND2_306 (N791, N708, N778);
nor NOR2_307 (N792, N717, N782);
and AND2_308 (N793, N717, N782);
and AND2_309 (N794, N219, N786);
  nand NAND2_310 (KeyWire_0[78], N628, N773);
  xor KeyGate_0_78(N795, keyIn_0_78, KeyWire_0[78]);
  nand NAND2_311 (KeyWire_0[79], N795, N747);
  xor KeyGate_0_79(KeyNOTWire_0[31], keyIn_0_79, KeyWire_0[79]);
  not KeyNOTGate_0_31(N796, KeyNOTWire_0[31]);
  nor NOR2_312 (KeyWire_0[80], N788, N789);
  xor KeyGate_0_80(KeyNOTWire_0[32], keyIn_0_80, KeyWire_0[80]);
  not KeyNOTGate_0_32(N802, KeyNOTWire_0[32]);
nor NOR2_313 (N803, N790, N791);
nor NOR2_314 (N804, N792, N793);
nor NOR2_315 (N805, N340, N794);
  nor NOR2_316 (KeyWire_0[81], N692, N796);
  xor KeyGate_0_81(KeyNOTWire_0[33], keyIn_0_81, KeyWire_0[81]);
  not KeyNOTGate_0_33(N806, KeyNOTWire_0[33]);
  and AND2_317 (KeyWire_0[82], N692, N796);
  xnor KeyGate_0_82(KeyNOTWire_0[34], keyIn_0_82, KeyWire_0[82]);
  not KeyNOTGate_0_34(N807, KeyNOTWire_0[34]);
  and AND2_318 (KeyWire_0[83], N219, N802);
  xor KeyGate_0_83(KeyNOTWire_0[35], keyIn_0_83, KeyWire_0[83]);
  not KeyNOTGate_0_35(N808, KeyNOTWire_0[35]);
and AND2_319 (N809, N219, N803);
  and AND2_320 (KeyWire_0[84], N219, N804);
  xor KeyGate_0_84(KeyNOTWire_0[36], keyIn_0_84, KeyWire_0[84]);
  not KeyNOTGate_0_36(N810, KeyNOTWire_0[36]);
nand NAND4_321 (N811, N805, N787, N731, N529);
  nand NAND2_322 (KeyWire_0[85], N619, N796);
  xor KeyGate_0_85(KeyNOTWire_0[37], keyIn_0_85, KeyWire_0[85]);
  not KeyNOTGate_0_37(N812, KeyNOTWire_0[37]);
  nand NAND3_323 (KeyWire_0[86], N609, N619, N796);
  xnor KeyGate_0_86(KeyNOTWire_0[38], keyIn_0_86, KeyWire_0[86]);
  not KeyNOTGate_0_38(N813, KeyNOTWire_0[38]);
  nand NAND4_324 (KeyWire_0[87], N600, N609, N619, N796);
  xnor KeyGate_0_87(KeyNOTWire_0[39], keyIn_0_87, KeyWire_0[87]);
  not KeyNOTGate_0_39(N814, KeyNOTWire_0[39]);
  nand NAND4_325 (KeyWire_0[88], N738, N765, N766, N814);
  xnor KeyGate_0_88(KeyNOTWire_0[40], keyIn_0_88, KeyWire_0[88]);
  not KeyNOTGate_0_40(N815, KeyNOTWire_0[40]);
  nand NAND3_326 (KeyWire_0[89], N741, N764, N813);
  xor KeyGate_0_89(KeyNOTWire_0[41], keyIn_0_89, KeyWire_0[89]);
  not KeyNOTGate_0_41(N819, KeyNOTWire_0[41]);
  nand NAND2_327 (KeyWire_0[90], N744, N812);
  xor KeyGate_0_90(N822, keyIn_0_90, KeyWire_0[90]);
  nor NOR2_328 (KeyWire_0[91], N806, N807);
  xnor KeyGate_0_91(KeyNOTWire_0[42], keyIn_0_91, KeyWire_0[91]);
  not KeyNOTGate_0_42(N825, KeyNOTWire_0[42]);
  nor NOR2_329 (KeyWire_0[92], N335, N808);
  xnor KeyGate_0_92(N826, keyIn_0_92, KeyWire_0[92]);
nor NOR2_330 (N827, N336, N809);
nor NOR2_331 (N828, N338, N810);
not NOT1_332 (N829, N811);
  nor NOR2_333 (KeyWire_0[93], N665, N815);
  xor KeyGate_0_93(KeyNOTWire_0[43], keyIn_0_93, KeyWire_0[93]);
  not KeyNOTGate_0_43(N830, KeyNOTWire_0[43]);
  and AND2_334 (KeyWire_0[94], N665, N815);
  xnor KeyGate_0_94(N831, keyIn_0_94, KeyWire_0[94]);
  nor NOR2_335 (KeyWire_0[95], N673, N819);
  xnor KeyGate_0_95(N832, keyIn_0_95, KeyWire_0[95]);
  and AND2_336 (KeyWire_0[96], N673, N819);
  xor KeyGate_0_96(N833, keyIn_0_96, KeyWire_0[96]);
  nor NOR2_337 (KeyWire_0[97], N682, N822);
  xor KeyGate_0_97(N834, keyIn_0_97, KeyWire_0[97]);
  and AND2_338 (KeyWire_0[98], N682, N822);
  xor KeyGate_0_98(N835, keyIn_0_98, KeyWire_0[98]);
  and AND2_339 (KeyWire_0[99], N219, N825);
  xnor KeyGate_0_99(N836, keyIn_0_99, KeyWire_0[99]);
  nand NAND3_340 (KeyWire_0[100], N826, N777, N704);
  xnor KeyGate_0_100(N837, keyIn_0_100, KeyWire_0[100]);
nand NAND4_341 (N838, N827, N781, N712, N527);
nand NAND4_342 (N839, N828, N785, N721, N528);
not NOT1_343 (N840, N829);
  nand NAND2_344 (KeyWire_0[101], N815, N593);
  xor KeyGate_0_101(KeyNOTWire_0[44], keyIn_0_101, KeyWire_0[101]);
  not KeyNOTGate_0_44(N841, KeyNOTWire_0[44]);
  nor NOR2_345 (KeyWire_0[102], N830, N831);
  xnor KeyGate_0_102(KeyNOTWire_0[45], keyIn_0_102, KeyWire_0[102]);
  not KeyNOTGate_0_45(N842, KeyNOTWire_0[45]);
  nor NOR2_346 (KeyWire_0[103], N832, N833);
  xnor KeyGate_0_103(N843, keyIn_0_103, KeyWire_0[103]);
  nor NOR2_347 (KeyWire_0[104], N834, N835);
  xor KeyGate_0_104(KeyNOTWire_0[46], keyIn_0_104, KeyWire_0[104]);
  not KeyNOTGate_0_46(N844, KeyNOTWire_0[46]);
  nor NOR2_348 (KeyWire_0[105], N334, N836);
  xor KeyGate_0_105(N845, keyIn_0_105, KeyWire_0[105]);
  not NOT1_349 (KeyWire_0[106], N837);
  xor KeyGate_0_106(KeyNOTWire_0[47], keyIn_0_106, KeyWire_0[106]);
  not KeyNOTGate_0_47(N846, KeyNOTWire_0[47]);
not NOT1_350 (N847, N838);
not NOT1_351 (N848, N839);
  and AND2_352 (KeyWire_0[107], N735, N841);
  xor KeyGate_0_107(N849, keyIn_0_107, KeyWire_0[107]);
buf BUFF1_353 (N850, N840);
  and AND2_354 (KeyWire_0[108], N219, N842);
  xnor KeyGate_0_108(N851, keyIn_0_108, KeyWire_0[108]);
  and AND2_355 (KeyWire_0[109], N219, N843);
  xnor KeyGate_0_109(N852, keyIn_0_109, KeyWire_0[109]);
  and AND2_356 (KeyWire_0[110], N219, N844);
  xor KeyGate_0_110(N853, keyIn_0_110, KeyWire_0[110]);
  nand NAND3_357 (KeyWire_0[111], N845, N772, N696);
  xnor KeyGate_0_111(N854, keyIn_0_111, KeyWire_0[111]);
  not NOT1_358 (KeyWire_0[112], N846);
  xor KeyGate_0_112(N855, keyIn_0_112, KeyWire_0[112]);
not NOT1_359 (N856, N847);
not NOT1_360 (N857, N848);
  not NOT1_361 (KeyWire_0[113], N849);
  xor KeyGate_0_113(KeyNOTWire_0[48], keyIn_0_113, KeyWire_0[113]);
  not KeyNOTGate_0_48(N858, KeyNOTWire_0[48]);
  nor NOR2_362 (KeyWire_0[114], N417, N851);
  xor KeyGate_0_114(N859, keyIn_0_114, KeyWire_0[114]);
  nor NOR2_363 (KeyWire_0[115], N332, N852);
  xor KeyGate_0_115(KeyNOTWire_0[49], keyIn_0_115, KeyWire_0[115]);
  not KeyNOTGate_0_49(N860, KeyNOTWire_0[49]);
  nor NOR2_364 (KeyWire_0[116], N333, N853);
  xor KeyGate_0_116(N861, keyIn_0_116, KeyWire_0[116]);
  not NOT1_365 (KeyWire_0[117], N854);
  xnor KeyGate_0_117(N862, keyIn_0_117, KeyWire_0[117]);
buf BUFF1_366 (N863, N855);
buf BUFF1_367 (N864, N856);
buf BUFF1_368 (N865, N857);
buf BUFF1_369 (N866, N858);
  nand NAND3_370 (KeyWire_0[118], N859, N769, N669);
  xnor KeyGate_0_118(N867, keyIn_0_118, KeyWire_0[118]);
  nand NAND3_371 (KeyWire_0[119], N860, N770, N677);
  xor KeyGate_0_119(KeyNOTWire_0[50], keyIn_0_119, KeyWire_0[119]);
  not KeyNOTGate_0_50(N868, KeyNOTWire_0[50]);
  nand NAND3_372 (KeyWire_0[120], N861, N771, N686);
  xnor KeyGate_0_120(KeyNOTWire_0[51], keyIn_0_120, KeyWire_0[120]);
  not KeyNOTGate_0_51(N869, KeyNOTWire_0[51]);
  not NOT1_373 (KeyWire_0[121], N862);
  xnor KeyGate_0_121(KeyNOTWire_0[52], keyIn_0_121, KeyWire_0[121]);
  not KeyNOTGate_0_52(N870, KeyNOTWire_0[52]);
  not NOT1_374 (KeyWire_0[122], N867);
  xor KeyGate_0_122(N871, keyIn_0_122, KeyWire_0[122]);
  not NOT1_375 (KeyWire_0[123], N868);
  xor KeyGate_0_123(N872, keyIn_0_123, KeyWire_0[123]);
  not NOT1_376 (KeyWire_0[124], N869);
  xnor KeyGate_0_124(N873, keyIn_0_124, KeyWire_0[124]);
buf BUFF1_377 (N874, N870);
  not NOT1_378 (KeyWire_0[125], N871);
  xor KeyGate_0_125(KeyNOTWire_0[53], keyIn_0_125, KeyWire_0[125]);
  not KeyNOTGate_0_53(N875, KeyNOTWire_0[53]);
  not NOT1_379 (KeyWire_0[126], N872);
  xnor KeyGate_0_126(N876, keyIn_0_126, KeyWire_0[126]);
  not NOT1_380 (KeyWire_0[127], N873);
  xor KeyGate_0_127(KeyNOTWire_0[54], keyIn_0_127, KeyWire_0[127]);
  not KeyNOTGate_0_54(N877, KeyNOTWire_0[54]);
buf BUFF1_381 (N878, N875);
buf BUFF1_382 (N879, N876);
buf BUFF1_383 (N880, N877);

endmodule
