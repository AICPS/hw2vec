`timescale 1ns / 1ps
// Verilog
// c1908
// Ninputs 33
// Noutputs 25
// NtotalGates 880
// NOT1 277
// NAND2 347
// BUFF1 162
// AND2 30
// AND3 12
// NAND4 2
// NAND3 1
// NAND8 3
// AND4 2
// NAND5 24
// AND5 16
// AND8 3
// NOR2 1

module top (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
                  N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899,
        keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4,
        keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9,
        keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14,
        keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19,
        keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24,
        keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29,
        keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34,
        keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39,
        keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44,
        keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49,
        keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54,
        keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59,
        keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64,
        keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69,
        keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74,
        keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79,
        keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84,
        keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89,
        keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94,
        keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99,
        keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104,
        keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109,
        keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114,
        keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119,
        keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124,
        keyIn_0_125, keyIn_0_126, keyIn_0_127);

  input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4;
  input keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9;
  input keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14;
  input keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19;
  input keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24;
  input keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29;
  input keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34;
  input keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39;
  input keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44;
  input keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49;
  input keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54;
  input keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59;
  input keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64;
  input keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69;
  input keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74;
  input keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79;
  input keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84;
  input keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89;
  input keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94;
  input keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99;
  input keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104;
  input keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109;
  input keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114;
  input keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119;
  input keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124;
  input keyIn_0_125, keyIn_0_126, keyIn_0_127;

  wire [0:127] KeyWire_0;
  wire [0:64] KeyNOTWire_0;

input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;

output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;

wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898;

not NOT1_1 (N190, N1);
not NOT1_2 (N194, N4);
not NOT1_3 (N197, N7);
  not NOT1_4 (KeyWire_0[0], N10);
  xor KeyGate_0_0(N201, keyIn_0_0, KeyWire_0[0]);
not NOT1_5 (N206, N13);
not NOT1_6 (N209, N16);
not NOT1_7 (N212, N19);
not NOT1_8 (N216, N22);
not NOT1_9 (N220, N25);
not NOT1_10 (N225, N28);
  not NOT1_11 (KeyWire_0[1], N31);
  xnor KeyGate_0_1(N229, keyIn_0_1, KeyWire_0[1]);
not NOT1_12 (N232, N34);
  not NOT1_13 (KeyWire_0[2], N37);
  xor KeyGate_0_2(KeyNOTWire_0[0], keyIn_0_2, KeyWire_0[2]);
  not KeyNOTGate_0_0(N235, KeyNOTWire_0[0]);
not NOT1_14 (N239, N40);
not NOT1_15 (N243, N43);
not NOT1_16 (N247, N46);
  nand NAND2_17 (KeyWire_0[3], N63, N88);
  xnor KeyGate_0_3(KeyNOTWire_0[1], keyIn_0_3, KeyWire_0[3]);
  not KeyNOTGate_0_1(N251, KeyNOTWire_0[1]);
nand NAND2_18 (N252, N66, N91);
not NOT1_19 (N253, N72);
not NOT1_20 (N256, N72);
buf BUFF1_21 (N257, N69);
buf BUFF1_22 (N260, N69);
not NOT1_23 (N263, N76);
not NOT1_24 (N266, N79);
not NOT1_25 (N269, N82);
  not NOT1_26 (KeyWire_0[4], N85);
  xor KeyGate_0_4(KeyNOTWire_0[2], keyIn_0_4, KeyWire_0[4]);
  not KeyNOTGate_0_2(N272, KeyNOTWire_0[2]);
not NOT1_27 (N275, N104);
not NOT1_28 (N276, N104);
not NOT1_29 (N277, N88);
not NOT1_30 (N280, N91);
buf BUFF1_31 (N283, N94);
not NOT1_32 (N290, N94);
buf BUFF1_33 (N297, N94);
not NOT1_34 (N300, N94);
buf BUFF1_35 (N303, N99);
not NOT1_36 (N306, N99);
not NOT1_37 (N313, N99);
buf BUFF1_38 (N316, N104);
not NOT1_39 (N319, N104);
buf BUFF1_40 (N326, N104);
buf BUFF1_41 (N331, N104);
not NOT1_42 (N338, N104);
buf BUFF1_43 (N343, N1);
buf BUFF1_44 (N346, N4);
buf BUFF1_45 (N349, N7);
buf BUFF1_46 (N352, N10);
buf BUFF1_47 (N355, N13);
buf BUFF1_48 (N358, N16);
buf BUFF1_49 (N361, N19);
buf BUFF1_50 (N364, N22);
buf BUFF1_51 (N367, N25);
buf BUFF1_52 (N370, N28);
buf BUFF1_53 (N373, N31);
buf BUFF1_54 (N376, N34);
buf BUFF1_55 (N379, N37);
buf BUFF1_56 (N382, N40);
buf BUFF1_57 (N385, N43);
buf BUFF1_58 (N388, N46);
not NOT1_59 (N534, N343);
not NOT1_60 (N535, N346);
not NOT1_61 (N536, N349);
not NOT1_62 (N537, N352);
not NOT1_63 (N538, N355);
not NOT1_64 (N539, N358);
not NOT1_65 (N540, N361);
not NOT1_66 (N541, N364);
not NOT1_67 (N542, N367);
not NOT1_68 (N543, N370);
not NOT1_69 (N544, N373);
not NOT1_70 (N545, N376);
not NOT1_71 (N546, N379);
not NOT1_72 (N547, N382);
not NOT1_73 (N548, N385);
not NOT1_74 (N549, N388);
  nand NAND2_75 (KeyWire_0[5], N306, N331);
  xnor KeyGate_0_5(N550, keyIn_0_5, KeyWire_0[5]);
nand NAND2_76 (N551, N306, N331);
  nand NAND2_77 (KeyWire_0[6], N306, N331);
  xnor KeyGate_0_6(KeyNOTWire_0[3], keyIn_0_6, KeyWire_0[6]);
  not KeyNOTGate_0_3(N552, KeyNOTWire_0[3]);
nand NAND2_78 (N553, N306, N331);
nand NAND2_79 (N554, N306, N331);
nand NAND2_80 (N555, N306, N331);
buf BUFF1_81 (N556, N190);
buf BUFF1_82 (N559, N194);
buf BUFF1_83 (N562, N206);
buf BUFF1_84 (N565, N209);
buf BUFF1_85 (N568, N225);
buf BUFF1_86 (N571, N243);
and AND2_87 (N574, N63, N319);
buf BUFF1_88 (N577, N220);
buf BUFF1_89 (N580, N229);
buf BUFF1_90 (N583, N232);
and AND2_91 (N586, N66, N319);
buf BUFF1_92 (N589, N239);
  and AND3_93 (KeyWire_0[7], N49, N253, N319);
  xnor KeyGate_0_7(N592, keyIn_0_7, KeyWire_0[7]);
buf BUFF1_94 (N595, N247);
buf BUFF1_95 (N598, N239);
nand NAND2_96 (N601, N326, N277);
nand NAND2_97 (N602, N326, N280);
nand NAND2_98 (N603, N260, N72);
nand NAND2_99 (N608, N260, N300);
nand NAND2_100 (N612, N256, N300);
buf BUFF1_101 (N616, N201);
buf BUFF1_102 (N619, N216);
buf BUFF1_103 (N622, N220);
buf BUFF1_104 (N625, N239);
buf BUFF1_105 (N628, N190);
buf BUFF1_106 (N631, N190);
buf BUFF1_107 (N634, N194);
buf BUFF1_108 (N637, N229);
buf BUFF1_109 (N640, N197);
and AND3_110 (N643, N56, N257, N319);
buf BUFF1_111 (N646, N232);
buf BUFF1_112 (N649, N201);
buf BUFF1_113 (N652, N235);
and AND3_114 (N655, N60, N257, N319);
buf BUFF1_115 (N658, N263);
buf BUFF1_116 (N661, N263);
buf BUFF1_117 (N664, N266);
buf BUFF1_118 (N667, N266);
buf BUFF1_119 (N670, N269);
buf BUFF1_120 (N673, N269);
buf BUFF1_121 (N676, N272);
buf BUFF1_122 (N679, N272);
and AND2_123 (N682, N251, N316);
and AND2_124 (N685, N252, N316);
buf BUFF1_125 (N688, N197);
buf BUFF1_126 (N691, N197);
buf BUFF1_127 (N694, N212);
buf BUFF1_128 (N697, N212);
buf BUFF1_129 (N700, N247);
buf BUFF1_130 (N703, N247);
buf BUFF1_131 (N706, N235);
buf BUFF1_132 (N709, N235);
buf BUFF1_133 (N712, N201);
buf BUFF1_134 (N715, N201);
buf BUFF1_135 (N718, N206);
buf BUFF1_136 (N721, N216);
and AND3_137 (N724, N53, N253, N319);
buf BUFF1_138 (N727, N243);
buf BUFF1_139 (N730, N220);
buf BUFF1_140 (N733, N220);
buf BUFF1_141 (N736, N209);
buf BUFF1_142 (N739, N216);
buf BUFF1_143 (N742, N225);
buf BUFF1_144 (N745, N243);
buf BUFF1_145 (N748, N212);
buf BUFF1_146 (N751, N225);
not NOT1_147 (N886, N682);
not NOT1_148 (N887, N685);
not NOT1_149 (N888, N616);
not NOT1_150 (N889, N619);
not NOT1_151 (N890, N622);
not NOT1_152 (N891, N625);
  not NOT1_153 (KeyWire_0[8], N631);
  xnor KeyGate_0_8(KeyNOTWire_0[4], keyIn_0_8, KeyWire_0[8]);
  not KeyNOTGate_0_4(N892, KeyNOTWire_0[4]);
not NOT1_154 (N893, N643);
not NOT1_155 (N894, N649);
  not NOT1_156 (KeyWire_0[9], N652);
  xor KeyGate_0_9(N895, keyIn_0_9, KeyWire_0[9]);
not NOT1_157 (N896, N655);
and AND2_158 (N897, N49, N612);
and AND2_159 (N898, N56, N608);
nand NAND2_160 (N899, N53, N612);
nand NAND2_161 (N903, N60, N608);
nand NAND2_162 (N907, N49, N612);
nand NAND2_163 (N910, N56, N608);
  not NOT1_164 (KeyWire_0[10], N661);
  xor KeyGate_0_10(KeyNOTWire_0[5], keyIn_0_10, KeyWire_0[10]);
  not KeyNOTGate_0_5(N913, KeyNOTWire_0[5]);
not NOT1_165 (N914, N658);
not NOT1_166 (N915, N667);
not NOT1_167 (N916, N664);
  not NOT1_168 (KeyWire_0[11], N673);
  xnor KeyGate_0_11(KeyNOTWire_0[6], keyIn_0_11, KeyWire_0[11]);
  not KeyNOTGate_0_6(N917, KeyNOTWire_0[6]);
not NOT1_169 (N918, N670);
  not NOT1_170 (KeyWire_0[12], N679);
  xnor KeyGate_0_12(KeyNOTWire_0[7], keyIn_0_12, KeyWire_0[12]);
  not KeyNOTGate_0_7(N919, KeyNOTWire_0[7]);
not NOT1_171 (N920, N676);
nand NAND4_172 (N921, N277, N297, N326, N603);
nand NAND4_173 (N922, N280, N297, N326, N603);
nand NAND3_174 (N923, N303, N338, N603);
and AND3_175 (N926, N303, N338, N603);
buf BUFF1_176 (N935, N556);
not NOT1_177 (N938, N688);
buf BUFF1_178 (N939, N556);
not NOT1_179 (N942, N691);
buf BUFF1_180 (N943, N562);
not NOT1_181 (N946, N694);
buf BUFF1_182 (N947, N562);
not NOT1_183 (N950, N697);
buf BUFF1_184 (N951, N568);
not NOT1_185 (N954, N700);
buf BUFF1_186 (N955, N568);
  not NOT1_187 (KeyWire_0[13], N703);
  xnor KeyGate_0_13(N958, keyIn_0_13, KeyWire_0[13]);
buf BUFF1_188 (N959, N574);
buf BUFF1_189 (N962, N574);
buf BUFF1_190 (N965, N580);
not NOT1_191 (N968, N706);
buf BUFF1_192 (N969, N580);
not NOT1_193 (N972, N709);
buf BUFF1_194 (N973, N586);
  not NOT1_195 (KeyWire_0[14], N712);
  xnor KeyGate_0_14(N976, keyIn_0_14, KeyWire_0[14]);
buf BUFF1_196 (N977, N586);
not NOT1_197 (N980, N715);
buf BUFF1_198 (N981, N592);
  not NOT1_199 (KeyWire_0[15], N628);
  xnor KeyGate_0_15(N984, keyIn_0_15, KeyWire_0[15]);
buf BUFF1_200 (N985, N592);
not NOT1_201 (N988, N718);
not NOT1_202 (N989, N721);
not NOT1_203 (N990, N634);
not NOT1_204 (N991, N724);
not NOT1_205 (N992, N727);
not NOT1_206 (N993, N637);
buf BUFF1_207 (N994, N595);
  not NOT1_208 (KeyWire_0[16], N730);
  xor KeyGate_0_16(N997, keyIn_0_16, KeyWire_0[16]);
buf BUFF1_209 (N998, N595);
not NOT1_210 (N1001, N733);
  not NOT1_211 (KeyWire_0[17], N736);
  xnor KeyGate_0_17(KeyNOTWire_0[8], keyIn_0_17, KeyWire_0[17]);
  not KeyNOTGate_0_8(N1002, KeyNOTWire_0[8]);
not NOT1_212 (N1003, N739);
not NOT1_213 (N1004, N640);
not NOT1_214 (N1005, N742);
not NOT1_215 (N1006, N745);
  not NOT1_216 (KeyWire_0[18], N646);
  xor KeyGate_0_18(N1007, keyIn_0_18, KeyWire_0[18]);
not NOT1_217 (N1008, N748);
not NOT1_218 (N1009, N751);
buf BUFF1_219 (N1010, N559);
buf BUFF1_220 (N1013, N559);
buf BUFF1_221 (N1016, N565);
buf BUFF1_222 (N1019, N565);
buf BUFF1_223 (N1022, N571);
buf BUFF1_224 (N1025, N571);
buf BUFF1_225 (N1028, N577);
buf BUFF1_226 (N1031, N577);
buf BUFF1_227 (N1034, N583);
buf BUFF1_228 (N1037, N583);
buf BUFF1_229 (N1040, N589);
buf BUFF1_230 (N1043, N589);
buf BUFF1_231 (N1046, N598);
buf BUFF1_232 (N1049, N598);
nand NAND2_233 (N1054, N619, N888);
nand NAND2_234 (N1055, N616, N889);
nand NAND2_235 (N1063, N625, N890);
nand NAND2_236 (N1064, N622, N891);
nand NAND2_237 (N1067, N655, N895);
nand NAND2_238 (N1068, N652, N896);
  nand NAND2_239 (KeyWire_0[19], N721, N988);
  xnor KeyGate_0_19(N1119, keyIn_0_19, KeyWire_0[19]);
nand NAND2_240 (N1120, N718, N989);
nand NAND2_241 (N1121, N727, N991);
nand NAND2_242 (N1122, N724, N992);
nand NAND2_243 (N1128, N739, N1002);
nand NAND2_244 (N1129, N736, N1003);
nand NAND2_245 (N1130, N745, N1005);
nand NAND2_246 (N1131, N742, N1006);
  nand NAND2_247 (KeyWire_0[20], N751, N1008);
  xnor KeyGate_0_20(N1132, keyIn_0_20, KeyWire_0[20]);
nand NAND2_248 (N1133, N748, N1009);
not NOT1_249 (N1148, N939);
  not NOT1_250 (KeyWire_0[21], N935);
  xor KeyGate_0_21(KeyNOTWire_0[9], keyIn_0_21, KeyWire_0[21]);
  not KeyNOTGate_0_9(N1149, KeyNOTWire_0[9]);
nand NAND2_251 (N1150, N1054, N1055);
not NOT1_252 (N1151, N943);
not NOT1_253 (N1152, N947);
not NOT1_254 (N1153, N955);
not NOT1_255 (N1154, N951);
not NOT1_256 (N1155, N962);
  not NOT1_257 (KeyWire_0[22], N969);
  xor KeyGate_0_22(N1156, keyIn_0_22, KeyWire_0[22]);
not NOT1_258 (N1157, N977);
nand NAND2_259 (N1158, N1063, N1064);
not NOT1_260 (N1159, N985);
nand NAND2_261 (N1160, N985, N892);
  not NOT1_262 (KeyWire_0[23], N998);
  xnor KeyGate_0_23(N1161, keyIn_0_23, KeyWire_0[23]);
nand NAND2_263 (N1162, N1067, N1068);
not NOT1_264 (N1163, N899);
buf BUFF1_265 (N1164, N899);
not NOT1_266 (N1167, N903);
buf BUFF1_267 (N1168, N903);
nand NAND2_268 (N1171, N921, N923);
nand NAND2_269 (N1188, N922, N923);
not NOT1_270 (N1205, N1010);
nand NAND2_271 (N1206, N1010, N938);
not NOT1_272 (N1207, N1013);
nand NAND2_273 (N1208, N1013, N942);
not NOT1_274 (N1209, N1016);
nand NAND2_275 (N1210, N1016, N946);
not NOT1_276 (N1211, N1019);
nand NAND2_277 (N1212, N1019, N950);
  not NOT1_278 (KeyWire_0[24], N1022);
  xor KeyGate_0_24(KeyNOTWire_0[10], keyIn_0_24, KeyWire_0[24]);
  not KeyNOTGate_0_10(N1213, KeyNOTWire_0[10]);
nand NAND2_279 (N1214, N1022, N954);
not NOT1_280 (N1215, N1025);
  nand NAND2_281 (KeyWire_0[25], N1025, N958);
  xnor KeyGate_0_25(N1216, keyIn_0_25, KeyWire_0[25]);
not NOT1_282 (N1217, N1028);
not NOT1_283 (N1218, N959);
not NOT1_284 (N1219, N1031);
not NOT1_285 (N1220, N1034);
nand NAND2_286 (N1221, N1034, N968);
not NOT1_287 (N1222, N965);
  not NOT1_288 (KeyWire_0[26], N1037);
  xnor KeyGate_0_26(N1223, keyIn_0_26, KeyWire_0[26]);
nand NAND2_289 (N1224, N1037, N972);
not NOT1_290 (N1225, N1040);
nand NAND2_291 (N1226, N1040, N976);
  not NOT1_292 (KeyWire_0[27], N973);
  xnor KeyGate_0_27(KeyNOTWire_0[11], keyIn_0_27, KeyWire_0[27]);
  not KeyNOTGate_0_11(N1227, KeyNOTWire_0[11]);
  not NOT1_293 (KeyWire_0[28], N1043);
  xnor KeyGate_0_28(N1228, keyIn_0_28, KeyWire_0[28]);
nand NAND2_294 (N1229, N1043, N980);
not NOT1_295 (N1230, N981);
nand NAND2_296 (N1231, N981, N984);
nand NAND2_297 (N1232, N1119, N1120);
nand NAND2_298 (N1235, N1121, N1122);
not NOT1_299 (N1238, N1046);
nand NAND2_300 (N1239, N1046, N997);
not NOT1_301 (N1240, N994);
not NOT1_302 (N1241, N1049);
nand NAND2_303 (N1242, N1049, N1001);
  nand NAND2_304 (KeyWire_0[29], N1128, N1129);
  xnor KeyGate_0_29(KeyNOTWire_0[12], keyIn_0_29, KeyWire_0[29]);
  not KeyNOTGate_0_12(N1243, KeyNOTWire_0[12]);
nand NAND2_305 (N1246, N1130, N1131);
nand NAND2_306 (N1249, N1132, N1133);
buf BUFF1_307 (N1252, N907);
buf BUFF1_308 (N1255, N907);
buf BUFF1_309 (N1258, N910);
buf BUFF1_310 (N1261, N910);
  not NOT1_311 (KeyWire_0[30], N1150);
  xnor KeyGate_0_30(N1264, keyIn_0_30, KeyWire_0[30]);
  nand NAND2_312 (KeyWire_0[31], N631, N1159);
  xor KeyGate_0_31(KeyNOTWire_0[13], keyIn_0_31, KeyWire_0[31]);
  not KeyNOTGate_0_13(N1267, KeyNOTWire_0[13]);
nand NAND2_313 (N1309, N688, N1205);
nand NAND2_314 (N1310, N691, N1207);
  nand NAND2_315 (KeyWire_0[32], N694, N1209);
  xnor KeyGate_0_32(N1311, keyIn_0_32, KeyWire_0[32]);
nand NAND2_316 (N1312, N697, N1211);
  nand NAND2_317 (KeyWire_0[33], N700, N1213);
  xnor KeyGate_0_33(KeyNOTWire_0[14], keyIn_0_33, KeyWire_0[33]);
  not KeyNOTGate_0_14(N1313, KeyNOTWire_0[14]);
nand NAND2_318 (N1314, N703, N1215);
nand NAND2_319 (N1315, N706, N1220);
nand NAND2_320 (N1316, N709, N1223);
nand NAND2_321 (N1317, N712, N1225);
nand NAND2_322 (N1318, N715, N1228);
not NOT1_323 (N1319, N1158);
nand NAND2_324 (N1322, N628, N1230);
nand NAND2_325 (N1327, N730, N1238);
nand NAND2_326 (N1328, N733, N1241);
  not NOT1_327 (KeyWire_0[34], N1162);
  xnor KeyGate_0_34(KeyNOTWire_0[15], keyIn_0_34, KeyWire_0[34]);
  not KeyNOTGate_0_15(N1334, KeyNOTWire_0[15]);
nand NAND2_328 (N1344, N1267, N1160);
nand NAND2_329 (N1345, N1249, N894);
not NOT1_330 (N1346, N1249);
  not NOT1_331 (KeyWire_0[35], N1255);
  xor KeyGate_0_35(N1348, keyIn_0_35, KeyWire_0[35]);
  not NOT1_332 (KeyWire_0[36], N1252);
  xor KeyGate_0_36(N1349, keyIn_0_36, KeyWire_0[36]);
not NOT1_333 (N1350, N1261);
  not NOT1_334 (KeyWire_0[37], N1258);
  xor KeyGate_0_37(N1351, keyIn_0_37, KeyWire_0[37]);
  nand NAND2_335 (KeyWire_0[38], N1309, N1206);
  xor KeyGate_0_38(KeyNOTWire_0[16], keyIn_0_38, KeyWire_0[38]);
  not KeyNOTGate_0_16(N1352, KeyNOTWire_0[16]);
  nand NAND2_336 (KeyWire_0[39], N1310, N1208);
  xnor KeyGate_0_39(N1355, keyIn_0_39, KeyWire_0[39]);
nand NAND2_337 (N1358, N1311, N1210);
nand NAND2_338 (N1361, N1312, N1212);
nand NAND2_339 (N1364, N1313, N1214);
nand NAND2_340 (N1367, N1314, N1216);
nand NAND2_341 (N1370, N1315, N1221);
nand NAND2_342 (N1373, N1316, N1224);
nand NAND2_343 (N1376, N1317, N1226);
nand NAND2_344 (N1379, N1318, N1229);
nand NAND2_345 (N1383, N1322, N1231);
not NOT1_346 (N1386, N1232);
nand NAND2_347 (N1387, N1232, N990);
not NOT1_348 (N1388, N1235);
nand NAND2_349 (N1389, N1235, N993);
nand NAND2_350 (N1390, N1327, N1239);
nand NAND2_351 (N1393, N1328, N1242);
not NOT1_352 (N1396, N1243);
  nand NAND2_353 (KeyWire_0[40], N1243, N1004);
  xor KeyGate_0_40(N1397, keyIn_0_40, KeyWire_0[40]);
not NOT1_354 (N1398, N1246);
nand NAND2_355 (N1399, N1246, N1007);
not NOT1_356 (N1409, N1319);
nand NAND2_357 (N1412, N649, N1346);
not NOT1_358 (N1413, N1334);
buf BUFF1_359 (N1416, N1264);
buf BUFF1_360 (N1419, N1264);
  nand NAND2_361 (KeyWire_0[41], N634, N1386);
  xnor KeyGate_0_41(KeyNOTWire_0[17], keyIn_0_41, KeyWire_0[41]);
  not KeyNOTGate_0_17(N1433, KeyNOTWire_0[17]);
nand NAND2_362 (N1434, N637, N1388);
nand NAND2_363 (N1438, N640, N1396);
  nand NAND2_364 (KeyWire_0[42], N646, N1398);
  xor KeyGate_0_42(KeyNOTWire_0[18], keyIn_0_42, KeyWire_0[42]);
  not KeyNOTGate_0_18(N1439, KeyNOTWire_0[18]);
  not NOT1_365 (KeyWire_0[43], N1344);
  xor KeyGate_0_43(N1440, keyIn_0_43, KeyWire_0[43]);
nand NAND2_366 (N1443, N1355, N1148);
not NOT1_367 (N1444, N1355);
  nand NAND2_368 (KeyWire_0[44], N1352, N1149);
  xnor KeyGate_0_44(KeyNOTWire_0[19], keyIn_0_44, KeyWire_0[44]);
  not KeyNOTGate_0_19(N1445, KeyNOTWire_0[19]);
  not NOT1_369 (KeyWire_0[45], N1352);
  xor KeyGate_0_45(N1446, keyIn_0_45, KeyWire_0[45]);
  nand NAND2_370 (KeyWire_0[46], N1358, N1151);
  xnor KeyGate_0_46(KeyNOTWire_0[20], keyIn_0_46, KeyWire_0[46]);
  not KeyNOTGate_0_20(N1447, KeyNOTWire_0[20]);
not NOT1_371 (N1448, N1358);
nand NAND2_372 (N1451, N1361, N1152);
not NOT1_373 (N1452, N1361);
nand NAND2_374 (N1453, N1367, N1153);
not NOT1_375 (N1454, N1367);
nand NAND2_376 (N1455, N1364, N1154);
not NOT1_377 (N1456, N1364);
  nand NAND2_378 (KeyWire_0[47], N1373, N1156);
  xnor KeyGate_0_47(N1457, keyIn_0_47, KeyWire_0[47]);
not NOT1_379 (N1458, N1373);
nand NAND2_380 (N1459, N1379, N1157);
not NOT1_381 (N1460, N1379);
  not NOT1_382 (KeyWire_0[48], N1383);
  xnor KeyGate_0_48(N1461, keyIn_0_48, KeyWire_0[48]);
nand NAND2_383 (N1462, N1393, N1161);
not NOT1_384 (N1463, N1393);
nand NAND2_385 (N1464, N1345, N1412);
not NOT1_386 (N1468, N1370);
nand NAND2_387 (N1469, N1370, N1222);
not NOT1_388 (N1470, N1376);
  nand NAND2_389 (KeyWire_0[49], N1376, N1227);
  xor KeyGate_0_49(KeyNOTWire_0[21], keyIn_0_49, KeyWire_0[49]);
  not KeyNOTGate_0_21(N1471, KeyNOTWire_0[21]);
nand NAND2_390 (N1472, N1387, N1433);
not NOT1_391 (N1475, N1390);
nand NAND2_392 (N1476, N1390, N1240);
nand NAND2_393 (N1478, N1389, N1434);
nand NAND2_394 (N1481, N1399, N1439);
nand NAND2_395 (N1484, N1397, N1438);
nand NAND2_396 (N1487, N939, N1444);
nand NAND2_397 (N1488, N935, N1446);
nand NAND2_398 (N1489, N943, N1448);
  not NOT1_399 (KeyWire_0[50], N1419);
  xnor KeyGate_0_50(N1490, keyIn_0_50, KeyWire_0[50]);
not NOT1_400 (N1491, N1416);
nand NAND2_401 (N1492, N947, N1452);
  nand NAND2_402 (KeyWire_0[51], N955, N1454);
  xnor KeyGate_0_51(N1493, keyIn_0_51, KeyWire_0[51]);
nand NAND2_403 (N1494, N951, N1456);
nand NAND2_404 (N1495, N969, N1458);
nand NAND2_405 (N1496, N977, N1460);
  nand NAND2_406 (KeyWire_0[52], N998, N1463);
  xor KeyGate_0_52(N1498, keyIn_0_52, KeyWire_0[52]);
  not NOT1_407 (KeyWire_0[53], N1440);
  xnor KeyGate_0_53(N1499, keyIn_0_53, KeyWire_0[53]);
nand NAND2_408 (N1500, N965, N1468);
  nand NAND2_409 (KeyWire_0[54], N973, N1470);
  xnor KeyGate_0_54(KeyNOTWire_0[22], keyIn_0_54, KeyWire_0[54]);
  not KeyNOTGate_0_22(N1501, KeyNOTWire_0[22]);
nand NAND2_410 (N1504, N994, N1475);
not NOT1_411 (N1510, N1464);
nand NAND2_412 (N1513, N1443, N1487);
nand NAND2_413 (N1514, N1445, N1488);
nand NAND2_414 (N1517, N1447, N1489);
nand NAND2_415 (N1520, N1451, N1492);
nand NAND2_416 (N1521, N1453, N1493);
  nand NAND2_417 (KeyWire_0[55], N1455, N1494);
  xor KeyGate_0_55(N1522, keyIn_0_55, KeyWire_0[55]);
nand NAND2_418 (N1526, N1457, N1495);
nand NAND2_419 (N1527, N1459, N1496);
not NOT1_420 (N1528, N1472);
nand NAND2_421 (N1529, N1462, N1498);
not NOT1_422 (N1530, N1478);
not NOT1_423 (N1531, N1481);
not NOT1_424 (N1532, N1484);
nand NAND2_425 (N1534, N1471, N1501);
nand NAND2_426 (N1537, N1469, N1500);
nand NAND2_427 (N1540, N1476, N1504);
not NOT1_428 (N1546, N1513);
  not NOT1_429 (KeyWire_0[56], N1521);
  xor KeyGate_0_56(KeyNOTWire_0[23], keyIn_0_56, KeyWire_0[56]);
  not KeyNOTGate_0_23(N1554, KeyNOTWire_0[23]);
not NOT1_430 (N1557, N1526);
not NOT1_431 (N1561, N1520);
  nand NAND2_432 (KeyWire_0[57], N1484, N1531);
  xor KeyGate_0_57(KeyNOTWire_0[24], keyIn_0_57, KeyWire_0[57]);
  not KeyNOTGate_0_24(N1567, KeyNOTWire_0[24]);
nand NAND2_433 (N1568, N1481, N1532);
not NOT1_434 (N1569, N1510);
not NOT1_435 (N1571, N1527);
not NOT1_436 (N1576, N1529);
buf BUFF1_437 (N1588, N1522);
not NOT1_438 (N1591, N1534);
not NOT1_439 (N1593, N1537);
nand NAND2_440 (N1594, N1540, N1530);
not NOT1_441 (N1595, N1540);
nand NAND2_442 (N1596, N1567, N1568);
buf BUFF1_443 (N1600, N1517);
buf BUFF1_444 (N1603, N1517);
buf BUFF1_445 (N1606, N1522);
buf BUFF1_446 (N1609, N1522);
buf BUFF1_447 (N1612, N1514);
buf BUFF1_448 (N1615, N1514);
buf BUFF1_449 (N1620, N1557);
buf BUFF1_450 (N1623, N1554);
not NOT1_451 (N1635, N1571);
nand NAND2_452 (N1636, N1478, N1595);
nand NAND2_453 (N1638, N1576, N1569);
  not NOT1_454 (KeyWire_0[58], N1576);
  xor KeyGate_0_58(KeyNOTWire_0[25], keyIn_0_58, KeyWire_0[58]);
  not KeyNOTGate_0_25(N1639, KeyNOTWire_0[25]);
buf BUFF1_455 (N1640, N1561);
buf BUFF1_456 (N1643, N1561);
buf BUFF1_457 (N1647, N1546);
buf BUFF1_458 (N1651, N1546);
buf BUFF1_459 (N1658, N1554);
buf BUFF1_460 (N1661, N1557);
buf BUFF1_461 (N1664, N1557);
nand NAND2_462 (N1671, N1596, N893);
not NOT1_463 (N1672, N1596);
not NOT1_464 (N1675, N1600);
not NOT1_465 (N1677, N1603);
nand NAND2_466 (N1678, N1606, N1217);
  not NOT1_467 (KeyWire_0[59], N1606);
  xnor KeyGate_0_59(N1679, keyIn_0_59, KeyWire_0[59]);
nand NAND2_468 (N1680, N1609, N1219);
not NOT1_469 (N1681, N1609);
not NOT1_470 (N1682, N1612);
not NOT1_471 (N1683, N1615);
nand NAND2_472 (N1685, N1594, N1636);
nand NAND2_473 (N1688, N1510, N1639);
buf BUFF1_474 (N1697, N1588);
buf BUFF1_475 (N1701, N1588);
nand NAND2_476 (N1706, N643, N1672);
not NOT1_477 (N1707, N1643);
nand NAND2_478 (N1708, N1647, N1675);
not NOT1_479 (N1709, N1647);
nand NAND2_480 (N1710, N1651, N1677);
  not NOT1_481 (KeyWire_0[60], N1651);
  xor KeyGate_0_60(N1711, keyIn_0_60, KeyWire_0[60]);
nand NAND2_482 (N1712, N1028, N1679);
nand NAND2_483 (N1713, N1031, N1681);
buf BUFF1_484 (N1714, N1620);
buf BUFF1_485 (N1717, N1620);
nand NAND2_486 (N1720, N1658, N1593);
not NOT1_487 (N1721, N1658);
nand NAND2_488 (N1723, N1638, N1688);
not NOT1_489 (N1727, N1661);
not NOT1_490 (N1728, N1640);
not NOT1_491 (N1730, N1664);
buf BUFF1_492 (N1731, N1623);
buf BUFF1_493 (N1734, N1623);
nand NAND2_494 (N1740, N1685, N1528);
  not NOT1_495 (KeyWire_0[61], N1685);
  xor KeyGate_0_61(KeyNOTWire_0[26], keyIn_0_61, KeyWire_0[61]);
  not KeyNOTGate_0_26(N1741, KeyNOTWire_0[26]);
nand NAND2_496 (N1742, N1671, N1706);
  nand NAND2_497 (KeyWire_0[62], N1600, N1709);
  xor KeyGate_0_62(KeyNOTWire_0[27], keyIn_0_62, KeyWire_0[62]);
  not KeyNOTGate_0_27(N1746, KeyNOTWire_0[27]);
nand NAND2_498 (N1747, N1603, N1711);
nand NAND2_499 (N1748, N1678, N1712);
nand NAND2_500 (N1751, N1680, N1713);
nand NAND2_501 (N1759, N1537, N1721);
not NOT1_502 (N1761, N1697);
nand NAND2_503 (N1762, N1697, N1727);
not NOT1_504 (N1763, N1701);
nand NAND2_505 (N1764, N1701, N1730);
not NOT1_506 (N1768, N1717);
nand NAND2_507 (N1769, N1472, N1741);
nand NAND2_508 (N1772, N1723, N1413);
not NOT1_509 (N1773, N1723);
  nand NAND2_510 (KeyWire_0[63], N1708, N1746);
  xor KeyGate_0_63(KeyNOTWire_0[28], keyIn_0_63, KeyWire_0[63]);
  not KeyNOTGate_0_28(N1774, KeyNOTWire_0[28]);
nand NAND2_511 (N1777, N1710, N1747);
not NOT1_512 (N1783, N1731);
nand NAND2_513 (N1784, N1731, N1682);
not NOT1_514 (N1785, N1714);
not NOT1_515 (N1786, N1734);
nand NAND2_516 (N1787, N1734, N1683);
nand NAND2_517 (N1788, N1720, N1759);
nand NAND2_518 (N1791, N1661, N1761);
nand NAND2_519 (N1792, N1664, N1763);
nand NAND2_520 (N1795, N1751, N1155);
not NOT1_521 (N1796, N1751);
  nand NAND2_522 (KeyWire_0[64], N1740, N1769);
  xor KeyGate_0_64(KeyNOTWire_0[29], keyIn_0_64, KeyWire_0[64]);
  not KeyNOTGate_0_29(N1798, KeyNOTWire_0[29]);
nand NAND2_523 (N1801, N1334, N1773);
nand NAND2_524 (N1802, N1742, N290);
not NOT1_525 (N1807, N1748);
nand NAND2_526 (N1808, N1748, N1218);
nand NAND2_527 (N1809, N1612, N1783);
nand NAND2_528 (N1810, N1615, N1786);
nand NAND2_529 (N1812, N1791, N1762);
nand NAND2_530 (N1815, N1792, N1764);
buf BUFF1_531 (N1818, N1742);
nand NAND2_532 (N1821, N1777, N1490);
not NOT1_533 (N1822, N1777);
nand NAND2_534 (N1823, N1774, N1491);
not NOT1_535 (N1824, N1774);
nand NAND2_536 (N1825, N962, N1796);
nand NAND2_537 (N1826, N1788, N1409);
not NOT1_538 (N1827, N1788);
  nand NAND2_539 (KeyWire_0[65], N1772, N1801);
  xor KeyGate_0_65(KeyNOTWire_0[30], keyIn_0_65, KeyWire_0[65]);
  not KeyNOTGate_0_30(N1830, KeyNOTWire_0[30]);
  nand NAND2_540 (KeyWire_0[66], N959, N1807);
  xnor KeyGate_0_66(N1837, keyIn_0_66, KeyWire_0[66]);
nand NAND2_541 (N1838, N1809, N1784);
nand NAND2_542 (N1841, N1810, N1787);
nand NAND2_543 (N1848, N1419, N1822);
nand NAND2_544 (N1849, N1416, N1824);
nand NAND2_545 (N1850, N1795, N1825);
  nand NAND2_546 (KeyWire_0[67], N1319, N1827);
  xnor KeyGate_0_67(KeyNOTWire_0[31], keyIn_0_67, KeyWire_0[67]);
  not KeyNOTGate_0_31(N1852, KeyNOTWire_0[31]);
nand NAND2_547 (N1855, N1815, N1707);
not NOT1_548 (N1856, N1815);
not NOT1_549 (N1857, N1818);
nand NAND2_550 (N1858, N1798, N290);
not NOT1_551 (N1864, N1812);
  nand NAND2_552 (KeyWire_0[68], N1812, N1728);
  xnor KeyGate_0_68(KeyNOTWire_0[32], keyIn_0_68, KeyWire_0[68]);
  not KeyNOTGate_0_32(N1865, KeyNOTWire_0[32]);
buf BUFF1_553 (N1866, N1798);
buf BUFF1_554 (N1869, N1802);
buf BUFF1_555 (N1872, N1802);
nand NAND2_556 (N1875, N1808, N1837);
nand NAND2_557 (N1878, N1821, N1848);
nand NAND2_558 (N1879, N1823, N1849);
nand NAND2_559 (N1882, N1841, N1768);
not NOT1_560 (N1883, N1841);
nand NAND2_561 (N1884, N1826, N1852);
  nand NAND2_562 (KeyWire_0[69], N1643, N1856);
  xnor KeyGate_0_69(KeyNOTWire_0[33], keyIn_0_69, KeyWire_0[69]);
  not KeyNOTGate_0_33(N1885, KeyNOTWire_0[33]);
nand NAND2_563 (N1889, N1830, N290);
not NOT1_564 (N1895, N1838);
nand NAND2_565 (N1896, N1838, N1785);
nand NAND2_566 (N1897, N1640, N1864);
  not NOT1_567 (KeyWire_0[70], N1850);
  xor KeyGate_0_70(KeyNOTWire_0[34], keyIn_0_70, KeyWire_0[70]);
  not KeyNOTGate_0_34(N1898, KeyNOTWire_0[34]);
buf BUFF1_568 (N1902, N1830);
not NOT1_569 (N1910, N1878);
  nand NAND2_570 (KeyWire_0[71], N1717, N1883);
  xnor KeyGate_0_71(KeyNOTWire_0[35], keyIn_0_71, KeyWire_0[71]);
  not KeyNOTGate_0_35(N1911, KeyNOTWire_0[35]);
  not NOT1_571 (KeyWire_0[72], N1884);
  xor KeyGate_0_72(KeyNOTWire_0[36], keyIn_0_72, KeyWire_0[72]);
  not KeyNOTGate_0_36(N1912, KeyNOTWire_0[36]);
  nand NAND2_572 (KeyWire_0[73], N1855, N1885);
  xor KeyGate_0_73(N1913, keyIn_0_73, KeyWire_0[73]);
not NOT1_573 (N1915, N1866);
nand NAND2_574 (N1919, N1872, N919);
not NOT1_575 (N1920, N1872);
  nand NAND2_576 (KeyWire_0[74], N1869, N920);
  xnor KeyGate_0_74(N1921, keyIn_0_74, KeyWire_0[74]);
not NOT1_577 (N1922, N1869);
not NOT1_578 (N1923, N1875);
nand NAND2_579 (N1924, N1714, N1895);
buf BUFF1_580 (N1927, N1858);
buf BUFF1_581 (N1930, N1858);
nand NAND2_582 (N1933, N1865, N1897);
nand NAND2_583 (N1936, N1882, N1911);
not NOT1_584 (N1937, N1898);
not NOT1_585 (N1938, N1902);
nand NAND2_586 (N1941, N679, N1920);
nand NAND2_587 (N1942, N676, N1922);
buf BUFF1_588 (N1944, N1879);
  not NOT1_589 (KeyWire_0[75], N1913);
  xor KeyGate_0_75(KeyNOTWire_0[37], keyIn_0_75, KeyWire_0[75]);
  not KeyNOTGate_0_37(N1947, KeyNOTWire_0[37]);
buf BUFF1_590 (N1950, N1889);
buf BUFF1_591 (N1953, N1889);
buf BUFF1_592 (N1958, N1879);
  nand NAND2_593 (KeyWire_0[76], N1896, N1924);
  xor KeyGate_0_76(KeyNOTWire_0[38], keyIn_0_76, KeyWire_0[76]);
  not KeyNOTGate_0_38(N1961, KeyNOTWire_0[38]);
and AND2_594 (N1965, N1910, N601);
and AND2_595 (N1968, N602, N1912);
nand NAND2_596 (N1975, N1930, N917);
not NOT1_597 (N1976, N1930);
nand NAND2_598 (N1977, N1927, N918);
not NOT1_599 (N1978, N1927);
nand NAND2_600 (N1979, N1919, N1941);
nand NAND2_601 (N1980, N1921, N1942);
not NOT1_602 (N1985, N1933);
not NOT1_603 (N1987, N1936);
not NOT1_604 (N1999, N1944);
nand NAND2_605 (N2000, N1944, N1937);
  not NOT1_606 (KeyWire_0[77], N1947);
  xnor KeyGate_0_77(KeyNOTWire_0[39], keyIn_0_77, KeyWire_0[77]);
  not KeyNOTGate_0_39(N2002, KeyNOTWire_0[39]);
nand NAND2_607 (N2003, N1947, N1499);
nand NAND2_608 (N2004, N1953, N1350);
not NOT1_609 (N2005, N1953);
nand NAND2_610 (N2006, N1950, N1351);
not NOT1_611 (N2007, N1950);
nand NAND2_612 (N2008, N673, N1976);
nand NAND2_613 (N2009, N670, N1978);
not NOT1_614 (N2012, N1979);
not NOT1_615 (N2013, N1958);
nand NAND2_616 (N2014, N1958, N1923);
not NOT1_617 (N2015, N1961);
nand NAND2_618 (N2016, N1961, N1635);
not NOT1_619 (N2018, N1965);
not NOT1_620 (N2019, N1968);
nand NAND2_621 (N2020, N1898, N1999);
  not NOT1_622 (KeyWire_0[78], N1987);
  xnor KeyGate_0_78(N2021, keyIn_0_78, KeyWire_0[78]);
nand NAND2_623 (N2022, N1987, N1591);
nand NAND2_624 (N2023, N1440, N2002);
nand NAND2_625 (N2024, N1261, N2005);
nand NAND2_626 (N2025, N1258, N2007);
nand NAND2_627 (N2026, N1975, N2008);
  nand NAND2_628 (KeyWire_0[79], N1977, N2009);
  xnor KeyGate_0_79(N2027, keyIn_0_79, KeyWire_0[79]);
not NOT1_629 (N2030, N1980);
buf BUFF1_630 (N2033, N1980);
nand NAND2_631 (N2036, N1875, N2013);
nand NAND2_632 (N2037, N1571, N2015);
nand NAND2_633 (N2038, N2020, N2000);
  nand NAND2_634 (KeyWire_0[80], N1534, N2021);
  xnor KeyGate_0_80(KeyNOTWire_0[40], keyIn_0_80, KeyWire_0[80]);
  not KeyNOTGate_0_40(N2039, KeyNOTWire_0[40]);
  nand NAND2_635 (KeyWire_0[81], N2023, N2003);
  xor KeyGate_0_81(KeyNOTWire_0[41], keyIn_0_81, KeyWire_0[81]);
  not KeyNOTGate_0_41(N2040, KeyNOTWire_0[41]);
  nand NAND2_636 (KeyWire_0[82], N2004, N2024);
  xor KeyGate_0_82(KeyNOTWire_0[42], keyIn_0_82, KeyWire_0[82]);
  not KeyNOTGate_0_42(N2041, KeyNOTWire_0[42]);
nand NAND2_637 (N2042, N2006, N2025);
not NOT1_638 (N2047, N2026);
nand NAND2_639 (N2052, N2036, N2014);
  nand NAND2_640 (KeyWire_0[83], N2037, N2016);
  xor KeyGate_0_83(KeyNOTWire_0[43], keyIn_0_83, KeyWire_0[83]);
  not KeyNOTGate_0_43(N2055, KeyNOTWire_0[43]);
not NOT1_641 (N2060, N2038);
nand NAND2_642 (N2061, N2039, N2022);
nand NAND2_643 (N2062, N2040, N290);
not NOT1_644 (N2067, N2041);
not NOT1_645 (N2068, N2027);
buf BUFF1_646 (N2071, N2027);
not NOT1_647 (N2076, N2052);
not NOT1_648 (N2077, N2055);
nand NAND2_649 (N2078, N2060, N290);
nand NAND2_650 (N2081, N2061, N290);
not NOT1_651 (N2086, N2042);
buf BUFF1_652 (N2089, N2042);
and AND2_653 (N2104, N2030, N2068);
  and AND2_654 (KeyWire_0[84], N2033, N2068);
  xor KeyGate_0_84(KeyNOTWire_0[44], keyIn_0_84, KeyWire_0[84]);
  not KeyNOTGate_0_44(N2119, KeyNOTWire_0[44]);
and AND2_655 (N2129, N2030, N2071);
and AND2_656 (N2143, N2033, N2071);
buf BUFF1_657 (N2148, N2062);
buf BUFF1_658 (N2151, N2062);
buf BUFF1_659 (N2196, N2078);
buf BUFF1_660 (N2199, N2078);
buf BUFF1_661 (N2202, N2081);
buf BUFF1_662 (N2205, N2081);
nand NAND2_663 (N2214, N2151, N915);
not NOT1_664 (N2215, N2151);
nand NAND2_665 (N2216, N2148, N916);
not NOT1_666 (N2217, N2148);
nand NAND2_667 (N2222, N2199, N1348);
not NOT1_668 (N2223, N2199);
nand NAND2_669 (N2224, N2196, N1349);
  not NOT1_670 (KeyWire_0[85], N2196);
  xor KeyGate_0_85(KeyNOTWire_0[45], keyIn_0_85, KeyWire_0[85]);
  not KeyNOTGate_0_45(N2225, KeyNOTWire_0[45]);
nand NAND2_671 (N2226, N2205, N913);
  not NOT1_672 (KeyWire_0[86], N2205);
  xnor KeyGate_0_86(KeyNOTWire_0[46], keyIn_0_86, KeyWire_0[86]);
  not KeyNOTGate_0_46(N2227, KeyNOTWire_0[46]);
  nand NAND2_673 (KeyWire_0[87], N2202, N914);
  xnor KeyGate_0_87(N2228, keyIn_0_87, KeyWire_0[87]);
not NOT1_674 (N2229, N2202);
nand NAND2_675 (N2230, N667, N2215);
nand NAND2_676 (N2231, N664, N2217);
nand NAND2_677 (N2232, N1255, N2223);
nand NAND2_678 (N2233, N1252, N2225);
nand NAND2_679 (N2234, N661, N2227);
nand NAND2_680 (N2235, N658, N2229);
nand NAND2_681 (N2236, N2214, N2230);
nand NAND2_682 (N2237, N2216, N2231);
nand NAND2_683 (N2240, N2222, N2232);
  nand NAND2_684 (KeyWire_0[88], N2224, N2233);
  xor KeyGate_0_88(KeyNOTWire_0[47], keyIn_0_88, KeyWire_0[88]);
  not KeyNOTGate_0_47(N2241, KeyNOTWire_0[47]);
nand NAND2_685 (N2244, N2226, N2234);
nand NAND2_686 (N2245, N2228, N2235);
not NOT1_687 (N2250, N2236);
  not NOT1_688 (KeyWire_0[89], N2240);
  xnor KeyGate_0_89(N2253, keyIn_0_89, KeyWire_0[89]);
not NOT1_689 (N2256, N2244);
not NOT1_690 (N2257, N2237);
buf BUFF1_691 (N2260, N2237);
  not NOT1_692 (KeyWire_0[90], N2241);
  xor KeyGate_0_90(N2263, keyIn_0_90, KeyWire_0[90]);
  and AND2_693 (KeyWire_0[91], N1164, N2241);
  xor KeyGate_0_91(KeyNOTWire_0[48], keyIn_0_91, KeyWire_0[91]);
  not KeyNOTGate_0_48(N2266, KeyNOTWire_0[48]);
not NOT1_694 (N2269, N2245);
and AND2_695 (N2272, N1168, N2245);
nand NAND8_696 (N2279, N2067, N2012, N2047, N2250, N899, N2256, N2253, N903);
buf BUFF1_697 (N2286, N2266);
buf BUFF1_698 (N2297, N2266);
buf BUFF1_699 (N2315, N2272);
buf BUFF1_700 (N2326, N2272);
and AND2_701 (N2340, N2086, N2257);
and AND2_702 (N2353, N2089, N2257);
  and AND2_703 (KeyWire_0[92], N2086, N2260);
  xnor KeyGate_0_92(N2361, keyIn_0_92, KeyWire_0[92]);
and AND2_704 (N2375, N2089, N2260);
  and AND4_705 (KeyWire_0[93], N338, N2279, N313, N313);
  xnor KeyGate_0_93(N2384, keyIn_0_93, KeyWire_0[93]);
and AND2_706 (N2385, N1163, N2263);
and AND2_707 (N2386, N1164, N2263);
and AND2_708 (N2426, N1167, N2269);
and AND2_709 (N2427, N1168, N2269);
nand NAND5_710 (N2537, N2286, N2315, N2361, N2104, N1171);
  nand NAND5_711 (KeyWire_0[94], N2286, N2315, N2340, N2129, N1171);
  xor KeyGate_0_94(N2540, keyIn_0_94, KeyWire_0[94]);
nand NAND5_712 (N2543, N2286, N2315, N2340, N2119, N1171);
nand NAND5_713 (N2546, N2286, N2315, N2353, N2104, N1171);
nand NAND5_714 (N2549, N2297, N2315, N2375, N2119, N1188);
nand NAND5_715 (N2552, N2297, N2326, N2361, N2143, N1188);
nand NAND5_716 (N2555, N2297, N2326, N2375, N2129, N1188);
and AND5_717 (N2558, N2286, N2315, N2361, N2104, N1171);
  and AND5_718 (KeyWire_0[95], N2286, N2315, N2340, N2129, N1171);
  xor KeyGate_0_95(KeyNOTWire_0[49], keyIn_0_95, KeyWire_0[95]);
  not KeyNOTGate_0_49(N2561, KeyNOTWire_0[49]);
and AND5_719 (N2564, N2286, N2315, N2340, N2119, N1171);
and AND5_720 (N2567, N2286, N2315, N2353, N2104, N1171);
and AND5_721 (N2570, N2297, N2315, N2375, N2119, N1188);
and AND5_722 (N2573, N2297, N2326, N2361, N2143, N1188);
  and AND5_723 (KeyWire_0[96], N2297, N2326, N2375, N2129, N1188);
  xnor KeyGate_0_96(KeyNOTWire_0[50], keyIn_0_96, KeyWire_0[96]);
  not KeyNOTGate_0_50(N2576, KeyNOTWire_0[50]);
nand NAND5_724 (N2594, N2286, N2427, N2361, N2129, N1171);
nand NAND5_725 (N2597, N2297, N2427, N2361, N2119, N1171);
nand NAND5_726 (N2600, N2297, N2427, N2375, N2104, N1171);
  nand NAND5_727 (KeyWire_0[97], N2297, N2427, N2340, N2143, N1171);
  xnor KeyGate_0_97(N2603, keyIn_0_97, KeyWire_0[97]);
  nand NAND5_728 (KeyWire_0[98], N2297, N2427, N2353, N2129, N1188);
  xor KeyGate_0_98(KeyNOTWire_0[51], keyIn_0_98, KeyWire_0[98]);
  not KeyNOTGate_0_51(N2606, KeyNOTWire_0[51]);
nand NAND5_729 (N2611, N2386, N2326, N2361, N2129, N1188);
nand NAND5_730 (N2614, N2386, N2326, N2361, N2119, N1188);
nand NAND5_731 (N2617, N2386, N2326, N2375, N2104, N1188);
nand NAND5_732 (N2620, N2386, N2326, N2353, N2129, N1188);
nand NAND5_733 (N2627, N2297, N2427, N2340, N2104, N926);
nand NAND5_734 (N2628, N2386, N2326, N2340, N2104, N926);
nand NAND5_735 (N2629, N2386, N2427, N2361, N2104, N926);
nand NAND5_736 (N2630, N2386, N2427, N2340, N2129, N926);
nand NAND5_737 (N2631, N2386, N2427, N2340, N2119, N926);
nand NAND5_738 (N2632, N2386, N2427, N2353, N2104, N926);
  nand NAND5_739 (KeyWire_0[99], N2386, N2426, N2340, N2104, N926);
  xor KeyGate_0_99(KeyNOTWire_0[52], keyIn_0_99, KeyWire_0[99]);
  not KeyNOTGate_0_52(N2633, KeyNOTWire_0[52]);
nand NAND5_740 (N2634, N2385, N2427, N2340, N2104, N926);
and AND5_741 (N2639, N2286, N2427, N2361, N2129, N1171);
  and AND5_742 (KeyWire_0[100], N2297, N2427, N2361, N2119, N1171);
  xnor KeyGate_0_100(KeyNOTWire_0[53], keyIn_0_100, KeyWire_0[100]);
  not KeyNOTGate_0_53(N2642, KeyNOTWire_0[53]);
and AND5_743 (N2645, N2297, N2427, N2375, N2104, N1171);
and AND5_744 (N2648, N2297, N2427, N2340, N2143, N1171);
and AND5_745 (N2651, N2297, N2427, N2353, N2129, N1188);
and AND5_746 (N2655, N2386, N2326, N2361, N2129, N1188);
  and AND5_747 (KeyWire_0[101], N2386, N2326, N2361, N2119, N1188);
  xnor KeyGate_0_101(N2658, keyIn_0_101, KeyWire_0[101]);
and AND5_748 (N2661, N2386, N2326, N2375, N2104, N1188);
  and AND5_749 (KeyWire_0[102], N2386, N2326, N2353, N2129, N1188);
  xnor KeyGate_0_102(N2664, keyIn_0_102, KeyWire_0[102]);
nand NAND2_750 (N2669, N2558, N534);
not NOT1_751 (N2670, N2558);
nand NAND2_752 (N2671, N2561, N535);
not NOT1_753 (N2672, N2561);
nand NAND2_754 (N2673, N2564, N536);
not NOT1_755 (N2674, N2564);
nand NAND2_756 (N2675, N2567, N537);
not NOT1_757 (N2676, N2567);
nand NAND2_758 (N2682, N2570, N543);
  not NOT1_759 (KeyWire_0[103], N2570);
  xnor KeyGate_0_103(KeyNOTWire_0[54], keyIn_0_103, KeyWire_0[103]);
  not KeyNOTGate_0_54(N2683, KeyNOTWire_0[54]);
nand NAND2_760 (N2688, N2573, N548);
  not NOT1_761 (KeyWire_0[104], N2573);
  xnor KeyGate_0_104(KeyNOTWire_0[55], keyIn_0_104, KeyWire_0[104]);
  not KeyNOTGate_0_55(N2689, KeyNOTWire_0[55]);
nand NAND2_762 (N2690, N2576, N549);
  not NOT1_763 (KeyWire_0[105], N2576);
  xor KeyGate_0_105(KeyNOTWire_0[56], keyIn_0_105, KeyWire_0[105]);
  not KeyNOTGate_0_56(N2691, KeyNOTWire_0[56]);
and AND8_764 (N2710, N2627, N2628, N2629, N2630, N2631, N2632, N2633, N2634);
nand NAND2_765 (N2720, N343, N2670);
nand NAND2_766 (N2721, N346, N2672);
nand NAND2_767 (N2722, N349, N2674);
nand NAND2_768 (N2723, N352, N2676);
  nand NAND2_769 (KeyWire_0[106], N2639, N538);
  xnor KeyGate_0_106(N2724, keyIn_0_106, KeyWire_0[106]);
not NOT1_770 (N2725, N2639);
  nand NAND2_771 (KeyWire_0[107], N2642, N539);
  xor KeyGate_0_107(KeyNOTWire_0[57], keyIn_0_107, KeyWire_0[107]);
  not KeyNOTGate_0_57(N2726, KeyNOTWire_0[57]);
not NOT1_772 (N2727, N2642);
nand NAND2_773 (N2728, N2645, N540);
not NOT1_774 (N2729, N2645);
nand NAND2_775 (N2730, N2648, N541);
not NOT1_776 (N2731, N2648);
nand NAND2_777 (N2732, N2651, N542);
  not NOT1_778 (KeyWire_0[108], N2651);
  xor KeyGate_0_108(KeyNOTWire_0[58], keyIn_0_108, KeyWire_0[108]);
  not KeyNOTGate_0_58(N2733, KeyNOTWire_0[58]);
  nand NAND2_779 (KeyWire_0[109], N370, N2683);
  xnor KeyGate_0_109(KeyNOTWire_0[59], keyIn_0_109, KeyWire_0[109]);
  not KeyNOTGate_0_59(N2734, KeyNOTWire_0[59]);
nand NAND2_780 (N2735, N2655, N544);
not NOT1_781 (N2736, N2655);
nand NAND2_782 (N2737, N2658, N545);
not NOT1_783 (N2738, N2658);
nand NAND2_784 (N2739, N2661, N546);
not NOT1_785 (N2740, N2661);
nand NAND2_786 (N2741, N2664, N547);
not NOT1_787 (N2742, N2664);
nand NAND2_788 (N2743, N385, N2689);
nand NAND2_789 (N2744, N388, N2691);
nand NAND8_790 (N2745, N2537, N2540, N2543, N2546, N2594, N2597, N2600, N2603);
nand NAND8_791 (N2746, N2606, N2549, N2611, N2614, N2617, N2620, N2552, N2555);
and AND8_792 (N2747, N2537, N2540, N2543, N2546, N2594, N2597, N2600, N2603);
and AND8_793 (N2750, N2606, N2549, N2611, N2614, N2617, N2620, N2552, N2555);
nand NAND2_794 (N2753, N2669, N2720);
nand NAND2_795 (N2754, N2671, N2721);
nand NAND2_796 (N2755, N2673, N2722);
  nand NAND2_797 (KeyWire_0[110], N2675, N2723);
  xnor KeyGate_0_110(N2756, keyIn_0_110, KeyWire_0[110]);
  nand NAND2_798 (KeyWire_0[111], N355, N2725);
  xor KeyGate_0_111(N2757, keyIn_0_111, KeyWire_0[111]);
  nand NAND2_799 (KeyWire_0[112], N358, N2727);
  xnor KeyGate_0_112(N2758, keyIn_0_112, KeyWire_0[112]);
nand NAND2_800 (N2759, N361, N2729);
nand NAND2_801 (N2760, N364, N2731);
nand NAND2_802 (N2761, N367, N2733);
nand NAND2_803 (N2762, N2682, N2734);
  nand NAND2_804 (KeyWire_0[113], N373, N2736);
  xor KeyGate_0_113(N2763, keyIn_0_113, KeyWire_0[113]);
nand NAND2_805 (N2764, N376, N2738);
nand NAND2_806 (N2765, N379, N2740);
nand NAND2_807 (N2766, N382, N2742);
  nand NAND2_808 (KeyWire_0[114], N2688, N2743);
  xnor KeyGate_0_114(N2767, keyIn_0_114, KeyWire_0[114]);
nand NAND2_809 (N2768, N2690, N2744);
and AND2_810 (N2773, N2745, N275);
and AND2_811 (N2776, N2746, N276);
  nand NAND2_812 (KeyWire_0[115], N2724, N2757);
  xor KeyGate_0_115(N2779, keyIn_0_115, KeyWire_0[115]);
nand NAND2_813 (N2780, N2726, N2758);
nand NAND2_814 (N2781, N2728, N2759);
nand NAND2_815 (N2782, N2730, N2760);
nand NAND2_816 (N2783, N2732, N2761);
nand NAND2_817 (N2784, N2735, N2763);
nand NAND2_818 (N2785, N2737, N2764);
  nand NAND2_819 (KeyWire_0[116], N2739, N2765);
  xor KeyGate_0_116(N2786, keyIn_0_116, KeyWire_0[116]);
nand NAND2_820 (N2787, N2741, N2766);
and AND3_821 (N2788, N2747, N2750, N2710);
nand NAND2_822 (N2789, N2747, N2750);
and AND4_823 (N2800, N338, N2279, N99, N2788);
  nand NAND2_824 (KeyWire_0[117], N2773, N2018);
  xor KeyGate_0_117(N2807, keyIn_0_117, KeyWire_0[117]);
not NOT1_825 (N2808, N2773);
  nand NAND2_826 (KeyWire_0[118], N2776, N2019);
  xnor KeyGate_0_118(N2809, keyIn_0_118, KeyWire_0[118]);
not NOT1_827 (N2810, N2776);
nor NOR2_828 (N2811, N2384, N2800);
and AND3_829 (N2812, N897, N283, N2789);
and AND3_830 (N2815, N76, N283, N2789);
  and AND3_831 (KeyWire_0[119], N82, N283, N2789);
  xor KeyGate_0_119(N2818, keyIn_0_119, KeyWire_0[119]);
and AND3_832 (N2821, N85, N283, N2789);
and AND3_833 (N2824, N898, N283, N2789);
nand NAND2_834 (N2827, N1965, N2808);
nand NAND2_835 (N2828, N1968, N2810);
  and AND3_836 (KeyWire_0[120], N79, N283, N2789);
  xnor KeyGate_0_120(N2829, keyIn_0_120, KeyWire_0[120]);
nand NAND2_837 (N2843, N2807, N2827);
nand NAND2_838 (N2846, N2809, N2828);
nand NAND2_839 (N2850, N2812, N2076);
nand NAND2_840 (N2851, N2815, N2077);
nand NAND2_841 (N2852, N2818, N1915);
  nand NAND2_842 (KeyWire_0[121], N2821, N1857);
  xor KeyGate_0_121(KeyNOTWire_0[60], keyIn_0_121, KeyWire_0[121]);
  not KeyNOTGate_0_60(N2853, KeyNOTWire_0[60]);
nand NAND2_843 (N2854, N2824, N1938);
not NOT1_844 (N2857, N2812);
  not NOT1_845 (KeyWire_0[122], N2815);
  xnor KeyGate_0_122(KeyNOTWire_0[61], keyIn_0_122, KeyWire_0[122]);
  not KeyNOTGate_0_61(N2858, KeyNOTWire_0[61]);
not NOT1_846 (N2859, N2818);
not NOT1_847 (N2860, N2821);
not NOT1_848 (N2861, N2824);
  not NOT1_849 (KeyWire_0[123], N2829);
  xnor KeyGate_0_123(N2862, keyIn_0_123, KeyWire_0[123]);
nand NAND2_850 (N2863, N2829, N1985);
nand NAND2_851 (N2866, N2052, N2857);
nand NAND2_852 (N2867, N2055, N2858);
  nand NAND2_853 (KeyWire_0[124], N1866, N2859);
  xnor KeyGate_0_124(KeyNOTWire_0[62], keyIn_0_124, KeyWire_0[124]);
  not KeyNOTGate_0_62(N2868, KeyNOTWire_0[62]);
nand NAND2_854 (N2869, N1818, N2860);
nand NAND2_855 (N2870, N1902, N2861);
nand NAND2_856 (N2871, N2843, N886);
  not NOT1_857 (KeyWire_0[125], N2843);
  xnor KeyGate_0_125(KeyNOTWire_0[63], keyIn_0_125, KeyWire_0[125]);
  not KeyNOTGate_0_63(N2872, KeyNOTWire_0[63]);
  nand NAND2_858 (KeyWire_0[126], N2846, N887);
  xnor KeyGate_0_126(N2873, keyIn_0_126, KeyWire_0[126]);
not NOT1_859 (N2874, N2846);
nand NAND2_860 (N2875, N1933, N2862);
nand NAND2_861 (N2876, N2866, N2850);
  nand NAND2_862 (KeyWire_0[127], N2867, N2851);
  xor KeyGate_0_127(KeyNOTWire_0[64], keyIn_0_127, KeyWire_0[127]);
  not KeyNOTGate_0_64(N2877, KeyNOTWire_0[64]);
nand NAND2_863 (N2878, N2868, N2852);
nand NAND2_864 (N2879, N2869, N2853);
nand NAND2_865 (N2880, N2870, N2854);
nand NAND2_866 (N2881, N682, N2872);
nand NAND2_867 (N2882, N685, N2874);
nand NAND2_868 (N2883, N2875, N2863);
and AND2_869 (N2886, N2876, N550);
and AND2_870 (N2887, N551, N2877);
and AND2_871 (N2888, N553, N2878);
and AND2_872 (N2889, N2879, N554);
and AND2_873 (N2890, N555, N2880);
nand NAND2_874 (N2891, N2871, N2881);
nand NAND2_875 (N2892, N2873, N2882);
nand NAND2_876 (N2895, N2883, N1461);
not NOT1_877 (N2896, N2883);
nand NAND2_878 (N2897, N1383, N2896);
nand NAND2_879 (N2898, N2895, N2897);
and AND2_880 (N2899, N2898, N552);

endmodule
