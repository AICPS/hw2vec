`timescale 1ns / 1ps
// Verilog
// c6288
// Ninputs 32
// Noutputs 32
// NtotalGates 2416
// AND2 256
// NOT1 32
// NOR2 2128

module top (N1,N18,N35,N52,N69,N86,N103,N120,N137,N154,
              N171,N188,N205,N222,N239,N256,N273,N290,N307,N324,
              N341,N358,N375,N392,N409,N426,N443,N460,N477,N494,
              N511,N528,N545,N1581,N1901,N2223,N2548,N2877,N3211,N3552,
              N3895,N4241,N4591,N4946,N5308,N5672,N5971,N6123,N6150,N6160,
              N6170,N6180,N6190,N6200,N6210,N6220,N6230,N6240,N6250,N6260,
                  N6270,N6280,N6287,N6288,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
        keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
        keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
        keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
        keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
        keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
        keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
        keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
        keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
        keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
        keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
        keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
        keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
        keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
        keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
        keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
        keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
        keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
                  keyinput255,
        keyinput256, keyinput257, keyinput258, keyinput259, keyinput260,
        keyinput261, keyinput262, keyinput263, keyinput264, keyinput265,
        keyinput266, keyinput267, keyinput268, keyinput269, keyinput270,
        keyinput271, keyinput272, keyinput273, keyinput274, keyinput275,
        keyinput276, keyinput277, keyinput278, keyinput279, keyinput280,
        keyinput281, keyinput282, keyinput283, keyinput284, keyinput285,
        keyinput286, keyinput287, keyinput288, keyinput289, keyinput290,
        keyinput291, keyinput292, keyinput293, keyinput294, keyinput295,
        keyinput296, keyinput297, keyinput298, keyinput299, keyinput300,
        keyinput301, keyinput302, keyinput303, keyinput304, keyinput305,
        keyinput306, keyinput307, keyinput308, keyinput309, keyinput310,
        keyinput311, keyinput312, keyinput313, keyinput314, keyinput315,
                  keyinput316, keyinput317, keyinput318, keyinput319,
        keyinput320, keyinput321, keyinput322, keyinput323, keyinput324,
        keyinput325, keyinput326, keyinput327, keyinput328, keyinput329,
        keyinput330, keyinput331, keyinput332, keyinput333, keyinput334,
        keyinput335, keyinput336, keyinput337, keyinput338, keyinput339,
        keyinput340, keyinput341, keyinput342, keyinput343, keyinput344,
        keyinput345, keyinput346, keyinput347, keyinput348, keyinput349,
        keyinput350, keyinput351);

  input keyinput320, keyinput321, keyinput322, keyinput323, keyinput324;
  input keyinput325, keyinput326, keyinput327, keyinput328, keyinput329;
  input keyinput330, keyinput331, keyinput332, keyinput333, keyinput334;
  input keyinput335, keyinput336, keyinput337, keyinput338, keyinput339;
  input keyinput340, keyinput341, keyinput342, keyinput343, keyinput344;
  input keyinput345, keyinput346, keyinput347, keyinput348, keyinput349;
  input keyinput350, keyinput351;


  input keyinput256, keyinput257, keyinput258, keyinput259, keyinput260;
  input keyinput261, keyinput262, keyinput263, keyinput264, keyinput265;
  input keyinput266, keyinput267, keyinput268, keyinput269, keyinput270;
  input keyinput271, keyinput272, keyinput273, keyinput274, keyinput275;
  input keyinput276, keyinput277, keyinput278, keyinput279, keyinput280;
  input keyinput281, keyinput282, keyinput283, keyinput284, keyinput285;
  input keyinput286, keyinput287, keyinput288, keyinput289, keyinput290;
  input keyinput291, keyinput292, keyinput293, keyinput294, keyinput295;
  input keyinput296, keyinput297, keyinput298, keyinput299, keyinput300;
  input keyinput301, keyinput302, keyinput303, keyinput304, keyinput305;
  input keyinput306, keyinput307, keyinput308, keyinput309, keyinput310;
  input keyinput311, keyinput312, keyinput313, keyinput314, keyinput315;
  input keyinput316, keyinput317, keyinput318, keyinput319;

  wire KeyWire_0_1 , KeyWire_0_2;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31, keyinput32, keyinput33, keyinput34;
  input keyinput35, keyinput36, keyinput37, keyinput38, keyinput39;
  input keyinput40, keyinput41, keyinput42, keyinput43, keyinput44;
  input keyinput45, keyinput46, keyinput47, keyinput48, keyinput49;
  input keyinput50, keyinput51, keyinput52, keyinput53, keyinput54;
  input keyinput55, keyinput56, keyinput57, keyinput58, keyinput59;
  input keyinput60, keyinput61, keyinput62, keyinput63, keyinput64;
  input keyinput65, keyinput66, keyinput67, keyinput68, keyinput69;
  input keyinput70, keyinput71, keyinput72, keyinput73, keyinput74;
  input keyinput75, keyinput76, keyinput77, keyinput78, keyinput79;
  input keyinput80, keyinput81, keyinput82, keyinput83, keyinput84;
  input keyinput85, keyinput86, keyinput87, keyinput88, keyinput89;
  input keyinput90, keyinput91, keyinput92, keyinput93, keyinput94;
  input keyinput95, keyinput96, keyinput97, keyinput98, keyinput99;
  input keyinput100, keyinput101, keyinput102, keyinput103, keyinput104;
  input keyinput105, keyinput106, keyinput107, keyinput108, keyinput109;
  input keyinput110, keyinput111, keyinput112, keyinput113, keyinput114;
  input keyinput115, keyinput116, keyinput117, keyinput118, keyinput119;
  input keyinput120, keyinput121, keyinput122, keyinput123, keyinput124;
  input keyinput125, keyinput126, keyinput127, keyinput128, keyinput129;
  input keyinput130, keyinput131, keyinput132, keyinput133, keyinput134;
  input keyinput135, keyinput136, keyinput137, keyinput138, keyinput139;
  input keyinput140, keyinput141, keyinput142, keyinput143, keyinput144;
  input keyinput145, keyinput146, keyinput147, keyinput148, keyinput149;
  input keyinput150, keyinput151, keyinput152, keyinput153, keyinput154;
  input keyinput155, keyinput156, keyinput157, keyinput158, keyinput159;
  input keyinput160, keyinput161, keyinput162, keyinput163, keyinput164;
  input keyinput165, keyinput166, keyinput167, keyinput168, keyinput169;
  input keyinput170, keyinput171, keyinput172, keyinput173, keyinput174;
  input keyinput175, keyinput176, keyinput177, keyinput178, keyinput179;
  input keyinput180, keyinput181, keyinput182, keyinput183, keyinput184;
  input keyinput185, keyinput186, keyinput187, keyinput188, keyinput189;
  input keyinput190, keyinput191, keyinput192, keyinput193, keyinput194;
  input keyinput195, keyinput196, keyinput197, keyinput198, keyinput199;
  input keyinput200, keyinput201, keyinput202, keyinput203, keyinput204;
  input keyinput205, keyinput206, keyinput207, keyinput208, keyinput209;
  input keyinput210, keyinput211, keyinput212, keyinput213, keyinput214;
  input keyinput215, keyinput216, keyinput217, keyinput218, keyinput219;
  input keyinput220, keyinput221, keyinput222, keyinput223, keyinput224;
  input keyinput225, keyinput226, keyinput227, keyinput228, keyinput229;
  input keyinput230, keyinput231, keyinput232, keyinput233, keyinput234;
  input keyinput235, keyinput236, keyinput237, keyinput238, keyinput239;
  input keyinput240, keyinput241, keyinput242, keyinput243, keyinput244;
  input keyinput245, keyinput246, keyinput247, keyinput248, keyinput249;
  input keyinput250, keyinput251, keyinput252, keyinput253, keyinput254;
  input keyinput255;

  wire [0:255] keyinput_Wire_0;
  wire [0:142] KeyNOTWire_0;

input N1,N18,N35,N52,N69,N86,N103,N120,N137,N154,
      N171,N188,N205,N222,N239,N256,N273,N290,N307,N324,
      N341,N358,N375,N392,N409,N426,N443,N460,N477,N494,
      N511,N528;

output N545,N1581,N1901,N2223,N2548,N2877,N3211,N3552,N3895,N4241,
       N4591,N4946,N5308,N5672,N5971,N6123,N6150,N6160,N6170,N6180,
       N6190,N6200,N6210,N6220,N6230,N6240,N6250,N6260,N6270,N6280,
       N6287,N6288;

wire N546,N549,N552,N555,N558,N561,N564,N567,N570,N573,
     N576,N579,N582,N585,N588,N591,N594,N597,N600,N603,
     N606,N609,N612,N615,N618,N621,N624,N627,N630,N633,
     N636,N639,N642,N645,N648,N651,N654,N657,N660,N663,
     N666,N669,N672,N675,N678,N681,N684,N687,N690,N693,
     N696,N699,N702,N705,N708,N711,N714,N717,N720,N723,
     N726,N729,N732,N735,N738,N741,N744,N747,N750,N753,
     N756,N759,N762,N765,N768,N771,N774,N777,N780,N783,
     N786,N789,N792,N795,N798,N801,N804,N807,N810,N813,
     N816,N819,N822,N825,N828,N831,N834,N837,N840,N843,
     N846,N849,N852,N855,N858,N861,N864,N867,N870,N873,
     N876,N879,N882,N885,N888,N891,N894,N897,N900,N903,
     N906,N909,N912,N915,N918,N921,N924,N927,N930,N933,
     N936,N939,N942,N945,N948,N951,N954,N957,N960,N963,
     N966,N969,N972,N975,N978,N981,N984,N987,N990,N993,
     N996,N999,N1002,N1005,N1008,N1011,N1014,N1017,N1020,N1023,
     N1026,N1029,N1032,N1035,N1038,N1041,N1044,N1047,N1050,N1053,
     N1056,N1059,N1062,N1065,N1068,N1071,N1074,N1077,N1080,N1083,
     N1086,N1089,N1092,N1095,N1098,N1101,N1104,N1107,N1110,N1113,
     N1116,N1119,N1122,N1125,N1128,N1131,N1134,N1137,N1140,N1143,
     N1146,N1149,N1152,N1155,N1158,N1161,N1164,N1167,N1170,N1173,
     N1176,N1179,N1182,N1185,N1188,N1191,N1194,N1197,N1200,N1203,
     N1206,N1209,N1212,N1215,N1218,N1221,N1224,N1227,N1230,N1233,
     N1236,N1239,N1242,N1245,N1248,N1251,N1254,N1257,N1260,N1263,
     N1266,N1269,N1272,N1275,N1278,N1281,N1284,N1287,N1290,N1293,
     N1296,N1299,N1302,N1305,N1308,N1311,N1315,N1319,N1323,N1327,
     N1331,N1335,N1339,N1343,N1347,N1351,N1355,N1359,N1363,N1367,
     N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,
     N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,
     N1391,N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,
     N1401,N1404,N1407,N1410,N1413,N1416,N1419,N1422,N1425,N1428,
     N1431,N1434,N1437,N1440,N1443,N1446,N1450,N1454,N1458,N1462,
     N1466,N1470,N1474,N1478,N1482,N1486,N1490,N1494,N1498,N1502,
     N1506,N1507,N1508,N1511,N1512,N1513,N1516,N1517,N1518,N1521,
     N1522,N1523,N1526,N1527,N1528,N1531,N1532,N1533,N1536,N1537,
     N1538,N1541,N1542,N1543,N1546,N1547,N1548,N1551,N1552,N1553,
     N1556,N1557,N1558,N1561,N1562,N1563,N1566,N1567,N1568,N1571,
     N1572,N1573,N1576,N1577,N1578,N1582,N1585,N1588,N1591,N1594,
     N1597,N1600,N1603,N1606,N1609,N1612,N1615,N1618,N1621,N1624,
     N1628,N1632,N1636,N1640,N1644,N1648,N1652,N1656,N1660,N1664,
     N1668,N1672,N1676,N1680,N1684,N1685,N1686,N1687,N1688,N1689,
     N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,
     N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,
     N1710,N1711,N1712,N1713,N1714,N1717,N1720,N1723,N1726,N1729,
     N1732,N1735,N1738,N1741,N1744,N1747,N1750,N1753,N1756,N1759,
     N1763,N1767,N1771,N1775,N1779,N1783,N1787,N1791,N1795,N1799,
     N1803,N1807,N1811,N1815,N1819,N1820,N1821,N1824,N1825,N1826,
     N1829,N1830,N1831,N1834,N1835,N1836,N1839,N1840,N1841,N1844,
     N1845,N1846,N1849,N1850,N1851,N1854,N1855,N1856,N1859,N1860,
     N1861,N1864,N1865,N1866,N1869,N1870,N1871,N1874,N1875,N1876,
     N1879,N1880,N1881,N1884,N1885,N1886,N1889,N1890,N1891,N1894,
     N1897,N1902,N1905,N1908,N1911,N1914,N1917,N1920,N1923,N1926,
     N1929,N1932,N1935,N1938,N1941,N1945,N1946,N1947,N1951,N1955,
     N1959,N1963,N1967,N1971,N1975,N1979,N1983,N1987,N1991,N1995,
     N1999,N2000,N2001,N2004,N2005,N2006,N2007,N2008,N2009,N2010,
     N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,
     N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,
     N2033,N2037,N2040,N2043,N2046,N2049,N2052,N2055,N2058,N2061,
     N2064,N2067,N2070,N2073,N2076,N2080,N2081,N2082,N2085,N2089,
     N2093,N2097,N2101,N2105,N2109,N2113,N2117,N2121,N2125,N2129,
     N2133,N2137,N2138,N2139,N2142,N2145,N2149,N2150,N2151,N2154,
     N2155,N2156,N2159,N2160,N2161,N2164,N2165,N2166,N2169,N2170,
     N2171,N2174,N2175,N2176,N2179,N2180,N2181,N2184,N2185,N2186,
     N2189,N2190,N2191,N2194,N2195,N2196,N2199,N2200,N2201,N2204,
     N2205,N2206,N2209,N2210,N2211,N2214,N2217,N2221,N2222,N2224,
     N2227,N2230,N2233,N2236,N2239,N2242,N2245,N2248,N2251,N2254,
     N2257,N2260,N2264,N2265,N2266,N2269,N2273,N2277,N2281,N2285,
     N2289,N2293,N2297,N2301,N2305,N2309,N2313,N2317,N2318,N2319,
     N2322,N2326,N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,
     N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,
     N2345,N2346,N2347,N2348,N2349,N2350,N2353,N2357,N2358,N2359,
     N2362,N2365,N2368,N2371,N2374,N2377,N2380,N2383,N2386,N2389,
     N2392,N2395,N2398,N2402,N2403,N2404,N2407,N2410,N2414,N2418,
     N2422,N2426,N2430,N2434,N2438,N2442,N2446,N2450,N2454,N2458,
     N2462,N2463,N2464,N2467,N2470,N2474,N2475,N2476,N2477,N2478,
     N2481,N2482,N2483,N2486,N2487,N2488,N2491,N2492,N2493,N2496,
     N2497,N2498,N2501,N2502,N2503,N2506,N2507,N2508,N2511,N2512,
     N2513,N2516,N2517,N2518,N2521,N2522,N2523,N2526,N2527,N2528,
     N2531,N2532,N2533,N2536,N2539,N2543,N2544,N2545,N2549,N2552,
     N2555,N2558,N2561,N2564,N2567,N2570,N2573,N2576,N2579,N2582,
     N2586,N2587,N2588,N2591,N2595,N2599,N2603,N2607,N2611,N2615,
     N2619,N2623,N2627,N2631,N2635,N2639,N2640,N2641,N2644,N2648,
     N2649,N2650,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,
     N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,
     N2671,N2672,N2673,N2674,N2675,N2678,N2682,N2683,N2684,N2687,
     N2690,N2694,N2697,N2700,N2703,N2706,N2709,N2712,N2715,N2718,
     N2721,N2724,N2727,N2731,N2732,N2733,N2736,N2739,N2743,N2744,
     N2745,N2749,N2753,N2757,N2761,N2765,N2769,N2773,N2777,N2781,
     N2785,N2789,N2790,N2791,N2794,N2797,N2801,N2802,N2803,N2806,
     N2807,N2808,N2811,N2812,N2813,N2816,N2817,N2818,N2821,N2822,
     N2823,N2826,N2827,N2828,N2831,N2832,N2833,N2836,N2837,N2838,
     N2841,N2842,N2843,N2846,N2847,N2848,N2851,N2852,N2853,N2856,
     N2857,N2858,N2861,N2864,N2868,N2869,N2870,N2873,N2878,N2881,
     N2884,N2887,N2890,N2893,N2896,N2899,N2902,N2905,N2908,N2912,
     N2913,N2914,N2917,N2921,N2922,N2923,N2926,N2930,N2934,N2938,
     N2942,N2946,N2950,N2954,N2958,N2962,N2966,N2967,N2968,N2971,
     N2975,N2976,N2977,N2980,N2983,N2987,N2988,N2989,N2990,N2991,
     N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,
     N3002,N3003,N3004,N3005,N3006,N3007,N3010,N3014,N3015,N3016,
     N3019,N3022,N3026,N3027,N3028,N3031,N3034,N3037,N3040,N3043,
     N3046,N3049,N3052,N3055,N3058,N3062,N3063,N3064,N3067,N3070,
     N3074,N3075,N3076,N3079,N3083,N3087,N3091,N3095,N3099,N3103,
     N3107,N3111,N3115,N3119,N3120,N3121,N3124,N3127,N3131,N3132,
     N3133,N3136,N3140,N3141,N3142,N3145,N3146,N3147,N3150,N3151,
     N3152,N3155,N3156,N3157,N3160,N3161,N3162,N3165,N3166,N3167,
     N3170,N3171,N3172,N3175,N3176,N3177,N3180,N3181,N3182,N3185,
     N3186,N3187,N3190,N3193,N3197,N3198,N3199,N3202,N3206,N3207,
     N3208,N3212,N3215,N3218,N3221,N3224,N3227,N3230,N3233,N3236,
     N3239,N3243,N3244,N3245,N3248,N3252,N3253,N3254,N3257,N3260,
     N3264,N3268,N3272,N3276,N3280,N3284,N3288,N3292,N3296,N3300,
     N3301,N3302,N3305,N3309,N3310,N3311,N3314,N3317,N3321,N3322,
     N3323,N3324,N3325,N3326,N3327,N3328,N3329,N3330,N3331,N3332,
     N3333,N3334,N3335,N3336,N3337,N3338,N3339,N3340,N3341,N3344,
     N3348,N3349,N3350,N3353,N3356,N3360,N3361,N3362,N3365,N3368,
     N3371,N3374,N3377,N3380,N3383,N3386,N3389,N3392,N3396,N3397,
     N3398,N3401,N3404,N3408,N3409,N3410,N3413,N3417,N3421,N3425,
     N3429,N3433,N3437,N3441,N3445,N3449,N3453,N3454,N3455,N3458,
     N3461,N3465,N3466,N3467,N3470,N3474,N3475,N3476,N3479,N3480,
     N3481,N3484,N3485,N3486,N3489,N3490,N3491,N3494,N3495,N3496,
     N3499,N3500,N3501,N3504,N3505,N3506,N3509,N3510,N3511,N3514,
     N3515,N3516,N3519,N3520,N3521,N3524,N3527,N3531,N3532,N3533,
     N3536,N3540,N3541,N3542,N3545,N3548,N3553,N3556,N3559,N3562,
     N3565,N3568,N3571,N3574,N3577,N3581,N3582,N3583,N3586,N3590,
     N3591,N3592,N3595,N3598,N3602,N3603,N3604,N3608,N3612,N3616,
     N3620,N3624,N3628,N3632,N3636,N3637,N3638,N3641,N3645,N3646,
     N3647,N3650,N3653,N3657,N3658,N3659,N3662,N3663,N3664,N3665,
     N3666,N3667,N3668,N3669,N3670,N3671,N3672,N3673,N3674,N3675,
     N3676,N3677,N3678,N3681,N3685,N3686,N3687,N3690,N3693,N3697,
     N3698,N3699,N3702,N3706,N3709,N3712,N3715,N3718,N3721,N3724,
     N3727,N3730,N3734,N3735,N3736,N3739,N3742,N3746,N3747,N3748,
     N3751,N3755,N3756,N3757,N3760,N3764,N3768,N3772,N3776,N3780,
     N3784,N3788,N3792,N3793,N3794,N3797,N3800,N3804,N3805,N3806,
     N3809,N3813,N3814,N3815,N3818,N3821,N3825,N3826,N3827,N3830,
     N3831,N3832,N3835,N3836,N3837,N3840,N3841,N3842,N3845,N3846,
     N3847,N3850,N3851,N3852,N3855,N3856,N3857,N3860,N3861,N3862,
     N3865,N3868,N3872,N3873,N3874,N3877,N3881,N3882,N3883,N3886,
     N3889,N3893,N3894,N3896,N3899,N3902,N3905,N3908,N3911,N3914,
     N3917,N3921,N3922,N3923,N3926,N3930,N3931,N3932,N3935,N3938,
     N3942,N3943,N3944,N3947,N3951,N3955,N3959,N3963,N3967,N3971,
     N3975,N3976,N3977,N3980,N3984,N3985,N3986,N3989,N3992,N3996,
     N3997,N3998,N4001,N4005,N4006,N4007,N4008,N4009,N4010,N4011,
     N4012,N4013,N4014,N4015,N4016,N4017,N4018,N4019,N4022,N4026,
     N4027,N4028,N4031,N4034,N4038,N4039,N4040,N4043,N4047,N4048,
     N4049,N4052,N4055,N4058,N4061,N4064,N4067,N4070,N4073,N4077,
     N4078,N4079,N4082,N4085,N4089,N4090,N4091,N4094,N4098,N4099,
     N4100,N4103,N4106,N4110,N4114,N4118,N4122,N4126,N4130,N4134,
     N4138,N4139,N4140,N4143,N4146,N4150,N4151,N4152,N4155,N4159,
     N4160,N4161,N4164,N4167,N4171,N4172,N4173,N4174,N4175,N4178,
     N4179,N4180,N4183,N4184,N4185,N4188,N4189,N4190,N4193,N4194,
     N4195,N4198,N4199,N4200,N4203,N4204,N4205,N4208,N4211,N4215,
     N4216,N4217,N4220,N4224,N4225,N4226,N4229,N4232,N4236,N4237,
     N4238,N4242,N4245,N4248,N4251,N4254,N4257,N4260,N4264,N4265,
     N4266,N4269,N4273,N4274,N4275,N4278,N4281,N4285,N4286,N4287,
     N4290,N4294,N4298,N4302,N4306,N4310,N4314,N4318,N4319,N4320,
     N4323,N4327,N4328,N4329,N4332,N4335,N4339,N4340,N4341,N4344,
     N4348,N4349,N4350,N4353,N4354,N4355,N4356,N4357,N4358,N4359,
     N4360,N4361,N4362,N4363,N4364,N4365,N4368,N4372,N4373,N4374,
     N4377,N4380,N4384,N4385,N4386,N4389,N4393,N4394,N4395,N4398,
     N4401,N4405,N4408,N4411,N4414,N4417,N4420,N4423,N4427,N4428,
     N4429,N4432,N4435,N4439,N4440,N4441,N4444,N4448,N4449,N4450,
     N4453,N4456,N4460,N4461,N4462,N4466,N4470,N4474,N4478,N4482,
     N4486,N4487,N4488,N4491,N4494,N4498,N4499,N4500,N4503,N4507,
     N4508,N4509,N4512,N4515,N4519,N4520,N4521,N4524,N4525,N4526,
     N4529,N4530,N4531,N4534,N4535,N4536,N4539,N4540,N4541,N4544,
     N4545,N4546,N4549,N4550,N4551,N4554,N4557,N4561,N4562,N4563,
     N4566,N4570,N4571,N4572,N4575,N4578,N4582,N4583,N4584,N4587,
     N4592,N4595,N4598,N4601,N4604,N4607,N4611,N4612,N4613,N4616,
     N4620,N4621,N4622,N4625,N4628,N4632,N4633,N4634,N4637,N4641,
     N4642,N4643,N4646,N4650,N4654,N4658,N4662,N4666,N4667,N4668,
     N4671,N4675,N4676,N4677,N4680,N4683,N4687,N4688,N4689,N4692,
     N4696,N4697,N4698,N4701,N4704,N4708,N4709,N4710,N4711,N4712,
     N4713,N4714,N4715,N4716,N4717,N4718,N4721,N4725,N4726,N4727,
     N4730,N4733,N4737,N4738,N4739,N4742,N4746,N4747,N4748,N4751,
     N4754,N4758,N4759,N4760,N4763,N4766,N4769,N4772,N4775,N4779,
     N4780,N4781,N4784,N4787,N4791,N4792,N4793,N4796,N4800,N4801,
     N4802,N4805,N4808,N4812,N4813,N4814,N4817,N4821,N4825,N4829,
     N4833,N4837,N4838,N4839,N4842,N4845,N4849,N4850,N4851,N4854,
     N4858,N4859,N4860,N4863,N4866,N4870,N4871,N4872,N4875,N4879,
     N4880,N4881,N4884,N4885,N4886,N4889,N4890,N4891,N4894,N4895,
     N4896,N4899,N4900,N4901,N4904,N4907,N4911,N4912,N4913,N4916,
     N4920,N4921,N4922,N4925,N4928,N4932,N4933,N4934,N4937,N4941,
     N4942,N4943,N4947,N4950,N4953,N4956,N4959,N4963,N4964,N4965,
     N4968,N4972,N4973,N4974,N4977,N4980,N4984,N4985,N4986,N4989,
     N4993,N4994,N4995,N4998,N5001,N5005,N5009,N5013,N5017,N5021,
     N5022,N5023,N5026,N5030,N5031,N5032,N5035,N5038,N5042,N5043,
     N5044,N5047,N5051,N5052,N5053,N5056,N5059,N5063,N5064,N5065,
     N5066,N5067,N5068,N5069,N5070,N5071,N5072,N5073,N5076,N5080,
     N5081,N5082,N5085,N5088,N5092,N5093,N5094,N5097,N5101,N5102,
     N5103,N5106,N5109,N5113,N5114,N5115,N5118,N5121,N5124,N5127,
     N5130,N5134,N5135,N5136,N5139,N5142,N5146,N5147,N5148,N5151,
     N5155,N5156,N5157,N5160,N5163,N5167,N5168,N5169,N5172,N5176,
     N5180,N5184,N5188,N5192,N5193,N5194,N5197,N5200,N5204,N5205,
     N5206,N5209,N5213,N5214,N5215,N5218,N5221,N5225,N5226,N5227,
     N5230,N5234,N5235,N5236,N5239,N5240,N5241,N5244,N5245,N5246,
     N5249,N5250,N5251,N5254,N5255,N5256,N5259,N5262,N5266,N5267,
     N5268,N5271,N5275,N5276,N5277,N5280,N5283,N5287,N5288,N5289,
     N5292,N5296,N5297,N5298,N5301,N5304,N5309,N5312,N5315,N5318,
     N5322,N5323,N5324,N5327,N5331,N5332,N5333,N5336,N5339,N5343,
     N5344,N5345,N5348,N5352,N5353,N5354,N5357,N5360,N5364,N5365,
     N5366,N5370,N5374,N5378,N5379,N5380,N5383,N5387,N5388,N5389,
     N5392,N5395,N5399,N5400,N5401,N5404,N5408,N5409,N5410,N5413,
     N5416,N5420,N5421,N5422,N5425,N5426,N5427,N5428,N5429,N5430,
     N5431,N5434,N5438,N5439,N5440,N5443,N5446,N5450,N5451,N5452,
     N5455,N5459,N5460,N5461,N5464,N5467,N5471,N5472,N5473,N5476,
     N5480,N5483,N5486,N5489,N5493,N5494,N5495,N5498,N5501,N5505,
     N5506,N5507,N5510,N5514,N5515,N5516,N5519,N5522,N5526,N5527,
     N5528,N5531,N5535,N5536,N5537,N5540,N5544,N5548,N5552,N5553,
     N5554,N5557,N5560,N5564,N5565,N5566,N5569,N5573,N5574,N5575,
     N5578,N5581,N5585,N5586,N5587,N5590,N5594,N5595,N5596,N5599,
     N5602,N5606,N5607,N5608,N5611,N5612,N5613,N5616,N5617,N5618,
     N5621,N5624,N5628,N5629,N5630,N5633,N5637,N5638,N5639,N5642,
     N5645,N5649,N5650,N5651,N5654,N5658,N5659,N5660,N5663,N5666,
     N5670,N5671,N5673,N5676,N5679,N5683,N5684,N5685,N5688,N5692,
     N5693,N5694,N5697,N5700,N5704,N5705,N5706,N5709,N5713,N5714,
     N5715,N5718,N5721,N5725,N5726,N5727,N5730,N5734,N5738,N5739,
     N5740,N5743,N5747,N5748,N5749,N5752,N5755,N5759,N5760,N5761,
     N5764,N5768,N5769,N5770,N5773,N5776,N5780,N5781,N5782,N5785,
     N5786,N5787,N5788,N5789,N5792,N5796,N5797,N5798,N5801,N5804,
     N5808,N5809,N5810,N5813,N5817,N5818,N5819,N5822,N5825,N5829,
     N5830,N5831,N5834,N5837,N5840,N5844,N5845,N5846,N5849,N5852,
     N5856,N5857,N5858,N5861,N5865,N5866,N5867,N5870,N5873,N5877,
     N5878,N5879,N5882,N5886,N5890,N5891,N5892,N5895,N5898,N5902,
     N5903,N5904,N5907,N5911,N5912,N5913,N5916,N5919,N5923,N5924,
     N5925,N5928,N5929,N5930,N5933,N5934,N5935,N5938,N5941,N5945,
     N5946,N5947,N5950,N5954,N5955,N5956,N5959,N5962,N5966,N5967,
     N5968,N5972,N5975,N5979,N5980,N5981,N5984,N5988,N5989,N5990,
     N5993,N5996,N6000,N6001,N6002,N6005,N6009,N6010,N6011,N6014,
     N6018,N6019,N6020,N6023,N6026,N6030,N6031,N6032,N6035,N6036,
     N6037,N6040,N6044,N6045,N6046,N6049,N6052,N6056,N6057,N6058,
     N6061,N6064,N6068,N6069,N6070,N6073,N6076,N6080,N6081,N6082,
     N6085,N6089,N6090,N6091,N6094,N6097,N6101,N6102,N6103,N6106,
     N6107,N6108,N6111,N6114,N6118,N6119,N6120,N6124,N6128,N6129,
     N6130,N6133,N6134,N6135,N6138,N6141,N6145,N6146,N6147,N6151,
     N6155,N6156,N6157,N6161,N6165,N6166,N6167,N6171,N6175,N6176,
     N6177,N6181,N6185,N6186,N6187,N6191,N6195,N6196,N6197,N6201,
     N6205,N6206,N6207,N6211,N6215,N6216,N6217,N6221,N6225,N6226,
     N6227,N6231,N6235,N6236,N6237,N6241,N6245,N6246,N6247,N6251,
     N6255,N6256,N6257,N6261,N6265,N6266,N6267,N6271,N6275,N6276,
     N6277,N6281,N6285,N6286;

and AND2_1 (N545, N1, N273);
and AND2_2 (N546, N1, N290);
and AND2_3 (N549, N1, N307);
and AND2_4 (N552, N1, N324);
and AND2_5 (N555, N1, N341);
and AND2_6 (N558, N1, N358);
and AND2_7 (N561, N1, N375);
and AND2_8 (N564, N1, N392);
and AND2_9 (N567, N1, N409);
and AND2_10 (N570, N1, N426);
and AND2_11 (N573, N1, N443);
and AND2_12 (N576, N1, N460);
and AND2_13 (N579, N1, N477);
and AND2_14 (N582, N1, N494);
and AND2_15 (N585, N1, N511);
and AND2_16 (N588, N1, N528);
and AND2_17 (N591, N18, N273);
and AND2_18 (N594, N18, N290);
and AND2_19 (N597, N18, N307);
and AND2_20 (N600, N18, N324);
and AND2_21 (N603, N18, N341);
and AND2_22 (N606, N18, N358);
and AND2_23 (N609, N18, N375);
and AND2_24 (N612, N18, N392);
and AND2_25 (N615, N18, N409);
and AND2_26 (N618, N18, N426);
and AND2_27 (N621, N18, N443);
and AND2_28 (N624, N18, N460);
and AND2_29 (N627, N18, N477);
and AND2_30 (N630, N18, N494);
and AND2_31 (N633, N18, N511);
and AND2_32 (N636, N18, N528);
and AND2_33 (N639, N35, N273);
and AND2_34 (N642, N35, N290);
and AND2_35 (N645, N35, N307);
and AND2_36 (N648, N35, N324);
and AND2_37 (N651, N35, N341);
and AND2_38 (N654, N35, N358);
and AND2_39 (N657, N35, N375);
and AND2_40 (N660, N35, N392);
and AND2_41 (N663, N35, N409);
and AND2_42 (N666, N35, N426);
and AND2_43 (N669, N35, N443);
and AND2_44 (N672, N35, N460);
and AND2_45 (N675, N35, N477);
and AND2_46 (N678, N35, N494);
and AND2_47 (N681, N35, N511);
and AND2_48 (N684, N35, N528);
and AND2_49 (N687, N52, N273);
and AND2_50 (N690, N52, N290);
and AND2_51 (N693, N52, N307);
and AND2_52 (N696, N52, N324);
and AND2_53 (N699, N52, N341);
and AND2_54 (N702, N52, N358);
and AND2_55 (N705, N52, N375);
and AND2_56 (N708, N52, N392);
and AND2_57 (N711, N52, N409);
and AND2_58 (N714, N52, N426);
and AND2_59 (N717, N52, N443);
and AND2_60 (N720, N52, N460);
and AND2_61 (N723, N52, N477);
and AND2_62 (N726, N52, N494);
and AND2_63 (N729, N52, N511);
and AND2_64 (N732, N52, N528);
and AND2_65 (N735, N69, N273);
and AND2_66 (N738, N69, N290);
and AND2_67 (N741, N69, N307);
and AND2_68 (N744, N69, N324);
and AND2_69 (N747, N69, N341);
and AND2_70 (N750, N69, N358);
and AND2_71 (N753, N69, N375);
and AND2_72 (N756, N69, N392);
and AND2_73 (N759, N69, N409);
and AND2_74 (N762, N69, N426);
and AND2_75 (N765, N69, N443);
and AND2_76 (N768, N69, N460);
and AND2_77 (N771, N69, N477);
and AND2_78 (N774, N69, N494);
and AND2_79 (N777, N69, N511);
and AND2_80 (N780, N69, N528);
and AND2_81 (N783, N86, N273);
and AND2_82 (N786, N86, N290);
and AND2_83 (N789, N86, N307);
and AND2_84 (N792, N86, N324);
and AND2_85 (N795, N86, N341);
and AND2_86 (N798, N86, N358);
and AND2_87 (N801, N86, N375);
and AND2_88 (N804, N86, N392);
and AND2_89 (N807, N86, N409);
and AND2_90 (N810, N86, N426);
and AND2_91 (N813, N86, N443);
and AND2_92 (N816, N86, N460);
and AND2_93 (N819, N86, N477);
and AND2_94 (N822, N86, N494);
and AND2_95 (N825, N86, N511);
  and AND2_96 (keyinput_Wire_0[0], N86, N528);
  xor keyGate_0_0(KeyNOTWire_0[0], keyinput0, keyinput_Wire_0[0]);
  not KeyNOTGate_0_0(N828, KeyNOTWire_0[0]);
and AND2_97 (N831, N103, N273);
and AND2_98 (N834, N103, N290);
and AND2_99 (N837, N103, N307);
and AND2_100 (N840, N103, N324);
and AND2_101 (N843, N103, N341);
and AND2_102 (N846, N103, N358);
and AND2_103 (N849, N103, N375);
and AND2_104 (N852, N103, N392);
and AND2_105 (N855, N103, N409);
and AND2_106 (N858, N103, N426);
and AND2_107 (N861, N103, N443);
and AND2_108 (N864, N103, N460);
and AND2_109 (N867, N103, N477);
and AND2_110 (N870, N103, N494);
and AND2_111 (N873, N103, N511);
and AND2_112 (N876, N103, N528);
and AND2_113 (N879, N120, N273);
and AND2_114 (N882, N120, N290);
and AND2_115 (N885, N120, N307);
and AND2_116 (N888, N120, N324);
and AND2_117 (N891, N120, N341);
and AND2_118 (N894, N120, N358);
and AND2_119 (N897, N120, N375);
and AND2_120 (N900, N120, N392);
and AND2_121 (N903, N120, N409);
and AND2_122 (N906, N120, N426);
and AND2_123 (N909, N120, N443);
and AND2_124 (N912, N120, N460);
and AND2_125 (N915, N120, N477);
and AND2_126 (N918, N120, N494);
and AND2_127 (N921, N120, N511);
and AND2_128 (N924, N120, N528);
and AND2_129 (N927, N137, N273);
and AND2_130 (N930, N137, N290);
and AND2_131 (N933, N137, N307);
and AND2_132 (N936, N137, N324);
and AND2_133 (N939, N137, N341);
and AND2_134 (N942, N137, N358);
and AND2_135 (N945, N137, N375);
and AND2_136 (N948, N137, N392);
and AND2_137 (N951, N137, N409);
and AND2_138 (N954, N137, N426);
and AND2_139 (N957, N137, N443);
and AND2_140 (N960, N137, N460);
and AND2_141 (N963, N137, N477);
and AND2_142 (N966, N137, N494);
and AND2_143 (N969, N137, N511);
and AND2_144 (N972, N137, N528);
and AND2_145 (N975, N154, N273);
and AND2_146 (N978, N154, N290);
and AND2_147 (N981, N154, N307);
and AND2_148 (N984, N154, N324);
and AND2_149 (N987, N154, N341);
and AND2_150 (N990, N154, N358);
and AND2_151 (N993, N154, N375);
and AND2_152 (N996, N154, N392);
and AND2_153 (N999, N154, N409);
and AND2_154 (N1002, N154, N426);
and AND2_155 (N1005, N154, N443);
and AND2_156 (N1008, N154, N460);
and AND2_157 (N1011, N154, N477);
and AND2_158 (N1014, N154, N494);
and AND2_159 (N1017, N154, N511);
and AND2_160 (N1020, N154, N528);
and AND2_161 (N1023, N171, N273);
  and AND2_162 (keyinput_Wire_0[1], N171, N290);
  xor keyGate_0_1(KeyNOTWire_0[1], keyinput1, keyinput_Wire_0[1]);
  not KeyNOTGate_0_1(N1026, KeyNOTWire_0[1]);
and AND2_163 (N1029, N171, N307);
and AND2_164 (N1032, N171, N324);
and AND2_165 (N1035, N171, N341);
and AND2_166 (N1038, N171, N358);
and AND2_167 (N1041, N171, N375);
and AND2_168 (N1044, N171, N392);
and AND2_169 (N1047, N171, N409);
and AND2_170 (N1050, N171, N426);
and AND2_171 (N1053, N171, N443);
and AND2_172 (N1056, N171, N460);
and AND2_173 (N1059, N171, N477);
and AND2_174 (N1062, N171, N494);
and AND2_175 (N1065, N171, N511);
and AND2_176 (N1068, N171, N528);
and AND2_177 (N1071, N188, N273);
and AND2_178 (N1074, N188, N290);
and AND2_179 (N1077, N188, N307);
and AND2_180 (N1080, N188, N324);
and AND2_181 (N1083, N188, N341);
and AND2_182 (N1086, N188, N358);
and AND2_183 (N1089, N188, N375);
and AND2_184 (N1092, N188, N392);
and AND2_185 (N1095, N188, N409);
and AND2_186 (N1098, N188, N426);
and AND2_187 (N1101, N188, N443);
and AND2_188 (N1104, N188, N460);
and AND2_189 (N1107, N188, N477);
and AND2_190 (N1110, N188, N494);
and AND2_191 (N1113, N188, N511);
and AND2_192 (N1116, N188, N528);
and AND2_193 (N1119, N205, N273);
and AND2_194 (N1122, N205, N290);
and AND2_195 (N1125, N205, N307);
and AND2_196 (N1128, N205, N324);
and AND2_197 (N1131, N205, N341);
and AND2_198 (N1134, N205, N358);
and AND2_199 (N1137, N205, N375);
and AND2_200 (N1140, N205, N392);
and AND2_201 (N1143, N205, N409);
and AND2_202 (N1146, N205, N426);
and AND2_203 (N1149, N205, N443);
and AND2_204 (N1152, N205, N460);
and AND2_205 (N1155, N205, N477);
and AND2_206 (N1158, N205, N494);
and AND2_207 (N1161, N205, N511);
and AND2_208 (N1164, N205, N528);
and AND2_209 (N1167, N222, N273);
  and AND2_210 (keyinput_Wire_0[2], N222, N290);
  xor keyGate_0_2(N1170, keyinput2, keyinput_Wire_0[2]);
  and AND2_211 (keyinput_Wire_0[3], N222, N307);
  xnor keyGate_0_3(N1173, keyinput3, keyinput_Wire_0[3]);
  and AND2_212 (keyinput_Wire_0[4], N222, N324);
  xor keyGate_0_4(KeyNOTWire_0[2], keyinput4, keyinput_Wire_0[4]);
  not KeyNOTGate_0_2(N1176, KeyNOTWire_0[2]);
  and AND2_213 (keyinput_Wire_0[5], N222, N341);
  xor keyGate_0_5(N1179, keyinput5, keyinput_Wire_0[5]);
  and AND2_214 (keyinput_Wire_0[6], N222, N358);
  xor keyGate_0_6(KeyNOTWire_0[3], keyinput6, keyinput_Wire_0[6]);
  not KeyNOTGate_0_3(N1182, KeyNOTWire_0[3]);
  and AND2_215 (keyinput_Wire_0[7], N222, N375);
  xor keyGate_0_7(N1185, keyinput7, keyinput_Wire_0[7]);
  and AND2_216 (keyinput_Wire_0[8], N222, N392);
  xor keyGate_0_8(N1188, keyinput8, keyinput_Wire_0[8]);
  and AND2_217 (keyinput_Wire_0[9], N222, N409);
  xor keyGate_0_9(N1191, keyinput9, keyinput_Wire_0[9]);
  and AND2_218 (keyinput_Wire_0[10], N222, N426);
  xnor keyGate_0_10(N1194, keyinput10, keyinput_Wire_0[10]);
  and AND2_219 (keyinput_Wire_0[11], N222, N443);
  xor keyGate_0_11(N1197, keyinput11, keyinput_Wire_0[11]);
  and AND2_220 (keyinput_Wire_0[12], N222, N460);
  xor keyGate_0_12(KeyNOTWire_0[4], keyinput12, keyinput_Wire_0[12]);
  not KeyNOTGate_0_4(N1200, KeyNOTWire_0[4]);
  and AND2_221 (keyinput_Wire_0[13], N222, N477);
  xor keyGate_0_13(KeyNOTWire_0[5], keyinput13, keyinput_Wire_0[13]);
  not KeyNOTGate_0_5(N1203, KeyNOTWire_0[5]);
  and AND2_222 (keyinput_Wire_0[14], N222, N494);
  xor keyGate_0_14(N1206, keyinput14, keyinput_Wire_0[14]);
and AND2_223 (N1209, N222, N511);
and AND2_224 (N1212, N222, N528);
  and AND2_225 (keyinput_Wire_0[15], N239, N273);
  xnor keyGate_0_15(N1215, keyinput15, keyinput_Wire_0[15]);
  and AND2_226 (keyinput_Wire_0[16], N239, N290);
  xnor keyGate_0_16(N1218, keyinput16, keyinput_Wire_0[16]);
  and AND2_227 (keyinput_Wire_0[17], N239, N307);
  xnor keyGate_0_17(N1221, keyinput17, keyinput_Wire_0[17]);
  and AND2_228 (keyinput_Wire_0[18], N239, N324);
  xor keyGate_0_18(N1224, keyinput18, keyinput_Wire_0[18]);
  and AND2_229 (keyinput_Wire_0[19], N239, N341);
  xor keyGate_0_19(KeyNOTWire_0[6], keyinput19, keyinput_Wire_0[19]);
  not KeyNOTGate_0_6(N1227, KeyNOTWire_0[6]);
  and AND2_230 (keyinput_Wire_0[20], N239, N358);
  xnor keyGate_0_20(N1230, keyinput20, keyinput_Wire_0[20]);
  and AND2_231 (keyinput_Wire_0[21], N239, N375);
  xor keyGate_0_21(KeyNOTWire_0[7], keyinput21, keyinput_Wire_0[21]);
  not KeyNOTGate_0_7(N1233, KeyNOTWire_0[7]);
  and AND2_232 (keyinput_Wire_0[22], N239, N392);
  xor keyGate_0_22(N1236, keyinput22, keyinput_Wire_0[22]);
  and AND2_233 (keyinput_Wire_0[23], N239, N409);
  xor keyGate_0_23(N1239, keyinput23, keyinput_Wire_0[23]);
  and AND2_234 (keyinput_Wire_0[24], N239, N426);
  xor keyGate_0_24(KeyNOTWire_0[8], keyinput24, keyinput_Wire_0[24]);
  not KeyNOTGate_0_8(N1242, KeyNOTWire_0[8]);
  and AND2_235 (keyinput_Wire_0[25], N239, N443);
  xor keyGate_0_25(KeyNOTWire_0[9], keyinput25, keyinput_Wire_0[25]);
  not KeyNOTGate_0_9(N1245, KeyNOTWire_0[9]);
  and AND2_236 (keyinput_Wire_0[26], N239, N460);
  xor keyGate_0_26(N1248, keyinput26, keyinput_Wire_0[26]);
  and AND2_237 (keyinput_Wire_0[27], N239, N477);
  xnor keyGate_0_27(KeyNOTWire_0[10], keyinput27, keyinput_Wire_0[27]);
  not KeyNOTGate_0_10(N1251, KeyNOTWire_0[10]);
  and AND2_238 (keyinput_Wire_0[28], N239, N494);
  xnor keyGate_0_28(KeyNOTWire_0[11], keyinput28, keyinput_Wire_0[28]);
  not KeyNOTGate_0_11(N1254, KeyNOTWire_0[11]);
and AND2_239 (N1257, N239, N511);
and AND2_240 (N1260, N239, N528);
  and AND2_241 (keyinput_Wire_0[29], N256, N273);
  xnor keyGate_0_29(KeyNOTWire_0[12], keyinput29, keyinput_Wire_0[29]);
  not KeyNOTGate_0_12(N1263, KeyNOTWire_0[12]);
  and AND2_242 (keyinput_Wire_0[30], N256, N290);
  xor keyGate_0_30(N1266, keyinput30, keyinput_Wire_0[30]);
  and AND2_243 (keyinput_Wire_0[31], N256, N307);
  xor keyGate_0_31(N1269, keyinput31, keyinput_Wire_0[31]);
  and AND2_244 (keyinput_Wire_0[32], N256, N324);
  xor keyGate_0_32(KeyNOTWire_0[13], keyinput32, keyinput_Wire_0[32]);
  not KeyNOTGate_0_13(N1272, KeyNOTWire_0[13]);
  and AND2_245 (keyinput_Wire_0[33], N256, N341);
  xnor keyGate_0_33(KeyNOTWire_0[14], keyinput33, keyinput_Wire_0[33]);
  not KeyNOTGate_0_14(N1275, KeyNOTWire_0[14]);
  and AND2_246 (keyinput_Wire_0[34], N256, N358);
  xnor keyGate_0_34(KeyNOTWire_0[15], keyinput34, keyinput_Wire_0[34]);
  not KeyNOTGate_0_15(N1278, KeyNOTWire_0[15]);
  and AND2_247 (keyinput_Wire_0[35], N256, N375);
  xor keyGate_0_35(KeyNOTWire_0[16], keyinput35, keyinput_Wire_0[35]);
  not KeyNOTGate_0_16(N1281, KeyNOTWire_0[16]);
  and AND2_248 (keyinput_Wire_0[36], N256, N392);
  xnor keyGate_0_36(KeyNOTWire_0[17], keyinput36, keyinput_Wire_0[36]);
  not KeyNOTGate_0_17(N1284, KeyNOTWire_0[17]);
  and AND2_249 (keyinput_Wire_0[37], N256, N409);
  xnor keyGate_0_37(N1287, keyinput37, keyinput_Wire_0[37]);
  and AND2_250 (keyinput_Wire_0[38], N256, N426);
  xnor keyGate_0_38(N1290, keyinput38, keyinput_Wire_0[38]);
  and AND2_251 (keyinput_Wire_0[39], N256, N443);
  xor keyGate_0_39(KeyNOTWire_0[18], keyinput39, keyinput_Wire_0[39]);
  not KeyNOTGate_0_18(N1293, KeyNOTWire_0[18]);
  and AND2_252 (keyinput_Wire_0[40], N256, N460);
  xnor keyGate_0_40(KeyNOTWire_0[19], keyinput40, keyinput_Wire_0[40]);
  not KeyNOTGate_0_19(N1296, KeyNOTWire_0[19]);
  and AND2_253 (keyinput_Wire_0[41], N256, N477);
  xnor keyGate_0_41(N1299, keyinput41, keyinput_Wire_0[41]);
and AND2_254 (N1302, N256, N494);
and AND2_255 (N1305, N256, N511);
and AND2_256 (N1308, N256, N528);
not NOT1_257 (N1311, N591);
  not NOT1_258 (keyinput_Wire_0[42], N639);
  xnor keyGate_0_42(N1315, keyinput42, keyinput_Wire_0[42]);
not NOT1_259 (N1319, N687);
not NOT1_260 (N1323, N735);
not NOT1_261 (N1327, N783);
not NOT1_262 (N1331, N831);
not NOT1_263 (N1335, N879);
not NOT1_264 (N1339, N927);
not NOT1_265 (N1343, N975);
not NOT1_266 (N1347, N1023);
not NOT1_267 (N1351, N1071);
not NOT1_268 (N1355, N1119);
not NOT1_269 (N1359, N1167);
  not NOT1_270 (keyinput_Wire_0[43], N1215);
  xor keyGate_0_43(KeyNOTWire_0[20], keyinput43, keyinput_Wire_0[43]);
  not KeyNOTGate_0_20(N1363, KeyNOTWire_0[20]);
  not NOT1_271 (keyinput_Wire_0[44], N1263);
  xnor keyGate_0_44(N1367, keyinput44, keyinput_Wire_0[44]);
nor NOR2_272 (N1371, N591, N1311);
not NOT1_273 (N1372, N1311);
nor NOR2_274 (N1373, N639, N1315);
not NOT1_275 (N1374, N1315);
nor NOR2_276 (N1375, N687, N1319);
not NOT1_277 (N1376, N1319);
nor NOR2_278 (N1377, N735, N1323);
not NOT1_279 (N1378, N1323);
nor NOR2_280 (N1379, N783, N1327);
not NOT1_281 (N1380, N1327);
nor NOR2_282 (N1381, N831, N1331);
not NOT1_283 (N1382, N1331);
nor NOR2_284 (N1383, N879, N1335);
not NOT1_285 (N1384, N1335);
nor NOR2_286 (N1385, N927, N1339);
not NOT1_287 (N1386, N1339);
nor NOR2_288 (N1387, N975, N1343);
not NOT1_289 (N1388, N1343);
nor NOR2_290 (N1389, N1023, N1347);
not NOT1_291 (N1390, N1347);
nor NOR2_292 (N1391, N1071, N1351);
not NOT1_293 (N1392, N1351);
nor NOR2_294 (N1393, N1119, N1355);
not NOT1_295 (N1394, N1355);
nor NOR2_296 (N1395, N1167, N1359);
not NOT1_297 (N1396, N1359);
  nor NOR2_298 (keyinput_Wire_0[45], N1215, N1363);
  xnor keyGate_0_45(KeyNOTWire_0[21], keyinput45, keyinput_Wire_0[45]);
  not KeyNOTGate_0_21(N1397, KeyNOTWire_0[21]);
  not NOT1_299 (keyinput_Wire_0[46], N1363);
  xor keyGate_0_46(N1398, keyinput46, keyinput_Wire_0[46]);
  nor NOR2_300 (keyinput_Wire_0[47], N1263, N1367);
  xnor keyGate_0_47(N1399, keyinput47, keyinput_Wire_0[47]);
  not NOT1_301 (keyinput_Wire_0[48], N1367);
  xnor keyGate_0_48(N1400, keyinput48, keyinput_Wire_0[48]);
nor NOR2_302 (N1401, N1371, N1372);
nor NOR2_303 (N1404, N1373, N1374);
nor NOR2_304 (N1407, N1375, N1376);
nor NOR2_305 (N1410, N1377, N1378);
nor NOR2_306 (N1413, N1379, N1380);
  nor NOR2_307 (keyinput_Wire_0[49], N1381, N1382);
  xor keyGate_0_49(KeyNOTWire_0[22], keyinput49, keyinput_Wire_0[49]);
  not KeyNOTGate_0_22(N1416, KeyNOTWire_0[22]);
nor NOR2_308 (N1419, N1383, N1384);
nor NOR2_309 (N1422, N1385, N1386);
nor NOR2_310 (N1425, N1387, N1388);
nor NOR2_311 (N1428, N1389, N1390);
nor NOR2_312 (N1431, N1391, N1392);
nor NOR2_313 (N1434, N1393, N1394);
nor NOR2_314 (N1437, N1395, N1396);
  nor NOR2_315 (keyinput_Wire_0[50], N1397, N1398);
  xor keyGate_0_50(KeyNOTWire_0[23], keyinput50, keyinput_Wire_0[50]);
  not KeyNOTGate_0_23(N1440, KeyNOTWire_0[23]);
  nor NOR2_316 (keyinput_Wire_0[51], N1399, N1400);
  xnor keyGate_0_51(N1443, keyinput51, keyinput_Wire_0[51]);
nor NOR2_317 (N1446, N1401, N546);
nor NOR2_318 (N1450, N1404, N594);
nor NOR2_319 (N1454, N1407, N642);
nor NOR2_320 (N1458, N1410, N690);
nor NOR2_321 (N1462, N1413, N738);
nor NOR2_322 (N1466, N1416, N786);
nor NOR2_323 (N1470, N1419, N834);
nor NOR2_324 (N1474, N1422, N882);
nor NOR2_325 (N1478, N1425, N930);
nor NOR2_326 (N1482, N1428, N978);
nor NOR2_327 (N1486, N1431, N1026);
nor NOR2_328 (N1490, N1434, N1074);
nor NOR2_329 (N1494, N1437, N1122);
  nor NOR2_330 (keyinput_Wire_0[52], N1440, N1170);
  xnor keyGate_0_52(N1498, keyinput52, keyinput_Wire_0[52]);
  nor NOR2_331 (keyinput_Wire_0[53], N1443, N1218);
  xor keyGate_0_53(KeyNOTWire_0[24], keyinput53, keyinput_Wire_0[53]);
  not KeyNOTGate_0_24(N1502, KeyNOTWire_0[24]);
nor NOR2_332 (N1506, N1401, N1446);
nor NOR2_333 (N1507, N1446, N546);
nor NOR2_334 (N1508, N1311, N1446);
nor NOR2_335 (N1511, N1404, N1450);
nor NOR2_336 (N1512, N1450, N594);
nor NOR2_337 (N1513, N1315, N1450);
nor NOR2_338 (N1516, N1407, N1454);
nor NOR2_339 (N1517, N1454, N642);
nor NOR2_340 (N1518, N1319, N1454);
nor NOR2_341 (N1521, N1410, N1458);
nor NOR2_342 (N1522, N1458, N690);
nor NOR2_343 (N1523, N1323, N1458);
nor NOR2_344 (N1526, N1413, N1462);
nor NOR2_345 (N1527, N1462, N738);
  nor NOR2_346 (keyinput_Wire_0[54], N1327, N1462);
  xnor keyGate_0_54(KeyNOTWire_0[25], keyinput54, keyinput_Wire_0[54]);
  not KeyNOTGate_0_25(N1528, KeyNOTWire_0[25]);
nor NOR2_347 (N1531, N1416, N1466);
nor NOR2_348 (N1532, N1466, N786);
nor NOR2_349 (N1533, N1331, N1466);
nor NOR2_350 (N1536, N1419, N1470);
nor NOR2_351 (N1537, N1470, N834);
nor NOR2_352 (N1538, N1335, N1470);
nor NOR2_353 (N1541, N1422, N1474);
nor NOR2_354 (N1542, N1474, N882);
nor NOR2_355 (N1543, N1339, N1474);
nor NOR2_356 (N1546, N1425, N1478);
nor NOR2_357 (N1547, N1478, N930);
nor NOR2_358 (N1548, N1343, N1478);
nor NOR2_359 (N1551, N1428, N1482);
nor NOR2_360 (N1552, N1482, N978);
nor NOR2_361 (N1553, N1347, N1482);
nor NOR2_362 (N1556, N1431, N1486);
nor NOR2_363 (N1557, N1486, N1026);
nor NOR2_364 (N1558, N1351, N1486);
nor NOR2_365 (N1561, N1434, N1490);
nor NOR2_366 (N1562, N1490, N1074);
nor NOR2_367 (N1563, N1355, N1490);
nor NOR2_368 (N1566, N1437, N1494);
nor NOR2_369 (N1567, N1494, N1122);
nor NOR2_370 (N1568, N1359, N1494);
nor NOR2_371 (N1571, N1440, N1498);
nor NOR2_372 (N1572, N1498, N1170);
  nor NOR2_373 (keyinput_Wire_0[55], N1363, N1498);
  xor keyGate_0_55(N1573, keyinput55, keyinput_Wire_0[55]);
  nor NOR2_374 (keyinput_Wire_0[56], N1443, N1502);
  xnor keyGate_0_56(KeyNOTWire_0[26], keyinput56, keyinput_Wire_0[56]);
  not KeyNOTGate_0_26(N1576, KeyNOTWire_0[26]);
  nor NOR2_375 (keyinput_Wire_0[57], N1502, N1218);
  xor keyGate_0_57(KeyNOTWire_0[27], keyinput57, keyinput_Wire_0[57]);
  not KeyNOTGate_0_27(N1577, KeyNOTWire_0[27]);
  nor NOR2_376 (keyinput_Wire_0[58], N1367, N1502);
  xor keyGate_0_58(KeyNOTWire_0[28], keyinput58, keyinput_Wire_0[58]);
  not KeyNOTGate_0_28(N1578, KeyNOTWire_0[28]);
nor NOR2_377 (N1581, N1506, N1507);
nor NOR2_378 (N1582, N1511, N1512);
nor NOR2_379 (N1585, N1516, N1517);
nor NOR2_380 (N1588, N1521, N1522);
nor NOR2_381 (N1591, N1526, N1527);
nor NOR2_382 (N1594, N1531, N1532);
nor NOR2_383 (N1597, N1536, N1537);
nor NOR2_384 (N1600, N1541, N1542);
nor NOR2_385 (N1603, N1546, N1547);
nor NOR2_386 (N1606, N1551, N1552);
nor NOR2_387 (N1609, N1556, N1557);
nor NOR2_388 (N1612, N1561, N1562);
nor NOR2_389 (N1615, N1566, N1567);
nor NOR2_390 (N1618, N1571, N1572);
  nor NOR2_391 (keyinput_Wire_0[59], N1576, N1577);
  xor keyGate_0_59(KeyNOTWire_0[29], keyinput59, keyinput_Wire_0[59]);
  not KeyNOTGate_0_29(N1621, KeyNOTWire_0[29]);
  nor NOR2_392 (keyinput_Wire_0[60], N1266, N1578);
  xor keyGate_0_60(KeyNOTWire_0[30], keyinput60, keyinput_Wire_0[60]);
  not KeyNOTGate_0_30(N1624, KeyNOTWire_0[30]);
nor NOR2_393 (N1628, N1582, N1508);
nor NOR2_394 (N1632, N1585, N1513);
nor NOR2_395 (N1636, N1588, N1518);
nor NOR2_396 (N1640, N1591, N1523);
nor NOR2_397 (N1644, N1594, N1528);
nor NOR2_398 (N1648, N1597, N1533);
nor NOR2_399 (N1652, N1600, N1538);
nor NOR2_400 (N1656, N1603, N1543);
  nor NOR2_401 (keyinput_Wire_0[61], N1606, N1548);
  xnor keyGate_0_61(N1660, keyinput61, keyinput_Wire_0[61]);
nor NOR2_402 (N1664, N1609, N1553);
nor NOR2_403 (N1668, N1612, N1558);
nor NOR2_404 (N1672, N1615, N1563);
nor NOR2_405 (N1676, N1618, N1568);
  nor NOR2_406 (keyinput_Wire_0[62], N1621, N1573);
  xor keyGate_0_62(KeyNOTWire_0[31], keyinput62, keyinput_Wire_0[62]);
  not KeyNOTGate_0_31(N1680, KeyNOTWire_0[31]);
  nor NOR2_407 (keyinput_Wire_0[63], N1266, N1624);
  xnor keyGate_0_63(KeyNOTWire_0[32], keyinput63, keyinput_Wire_0[63]);
  not KeyNOTGate_0_32(N1684, KeyNOTWire_0[32]);
  nor NOR2_408 (keyinput_Wire_0[64], N1624, N1578);
  xnor keyGate_0_64(KeyNOTWire_0[33], keyinput64, keyinput_Wire_0[64]);
  not KeyNOTGate_0_33(N1685, KeyNOTWire_0[33]);
nor NOR2_409 (N1686, N1582, N1628);
nor NOR2_410 (N1687, N1628, N1508);
nor NOR2_411 (N1688, N1585, N1632);
nor NOR2_412 (N1689, N1632, N1513);
nor NOR2_413 (N1690, N1588, N1636);
nor NOR2_414 (N1691, N1636, N1518);
nor NOR2_415 (N1692, N1591, N1640);
nor NOR2_416 (N1693, N1640, N1523);
nor NOR2_417 (N1694, N1594, N1644);
nor NOR2_418 (N1695, N1644, N1528);
nor NOR2_419 (N1696, N1597, N1648);
nor NOR2_420 (N1697, N1648, N1533);
nor NOR2_421 (N1698, N1600, N1652);
nor NOR2_422 (N1699, N1652, N1538);
nor NOR2_423 (N1700, N1603, N1656);
nor NOR2_424 (N1701, N1656, N1543);
nor NOR2_425 (N1702, N1606, N1660);
  nor NOR2_426 (keyinput_Wire_0[65], N1660, N1548);
  xor keyGate_0_65(N1703, keyinput65, keyinput_Wire_0[65]);
nor NOR2_427 (N1704, N1609, N1664);
nor NOR2_428 (N1705, N1664, N1553);
nor NOR2_429 (N1706, N1612, N1668);
nor NOR2_430 (N1707, N1668, N1558);
nor NOR2_431 (N1708, N1615, N1672);
nor NOR2_432 (N1709, N1672, N1563);
nor NOR2_433 (N1710, N1618, N1676);
nor NOR2_434 (N1711, N1676, N1568);
  nor NOR2_435 (keyinput_Wire_0[66], N1621, N1680);
  xor keyGate_0_66(N1712, keyinput66, keyinput_Wire_0[66]);
  nor NOR2_436 (keyinput_Wire_0[67], N1680, N1573);
  xor keyGate_0_67(N1713, keyinput67, keyinput_Wire_0[67]);
  nor NOR2_437 (keyinput_Wire_0[68], N1684, N1685);
  xor keyGate_0_68(N1714, keyinput68, keyinput_Wire_0[68]);
nor NOR2_438 (N1717, N1686, N1687);
nor NOR2_439 (N1720, N1688, N1689);
nor NOR2_440 (N1723, N1690, N1691);
nor NOR2_441 (N1726, N1692, N1693);
nor NOR2_442 (N1729, N1694, N1695);
nor NOR2_443 (N1732, N1696, N1697);
nor NOR2_444 (N1735, N1698, N1699);
nor NOR2_445 (N1738, N1700, N1701);
nor NOR2_446 (N1741, N1702, N1703);
nor NOR2_447 (N1744, N1704, N1705);
nor NOR2_448 (N1747, N1706, N1707);
nor NOR2_449 (N1750, N1708, N1709);
nor NOR2_450 (N1753, N1710, N1711);
  nor NOR2_451 (keyinput_Wire_0[69], N1712, N1713);
  xor keyGate_0_69(KeyNOTWire_0[34], keyinput69, keyinput_Wire_0[69]);
  not KeyNOTGate_0_34(N1756, KeyNOTWire_0[34]);
  nor NOR2_452 (keyinput_Wire_0[70], N1714, N1221);
  xor keyGate_0_70(KeyNOTWire_0[35], keyinput70, keyinput_Wire_0[70]);
  not KeyNOTGate_0_35(N1759, KeyNOTWire_0[35]);
nor NOR2_453 (N1763, N1717, N549);
nor NOR2_454 (N1767, N1720, N597);
nor NOR2_455 (N1771, N1723, N645);
nor NOR2_456 (N1775, N1726, N693);
nor NOR2_457 (N1779, N1729, N741);
nor NOR2_458 (N1783, N1732, N789);
  nor NOR2_459 (keyinput_Wire_0[71], N1735, N837);
  xor keyGate_0_71(KeyNOTWire_0[36], keyinput71, keyinput_Wire_0[71]);
  not KeyNOTGate_0_36(N1787, KeyNOTWire_0[36]);
nor NOR2_460 (N1791, N1738, N885);
nor NOR2_461 (N1795, N1741, N933);
nor NOR2_462 (N1799, N1744, N981);
nor NOR2_463 (N1803, N1747, N1029);
nor NOR2_464 (N1807, N1750, N1077);
nor NOR2_465 (N1811, N1753, N1125);
  nor NOR2_466 (keyinput_Wire_0[72], N1756, N1173);
  xnor keyGate_0_72(KeyNOTWire_0[37], keyinput72, keyinput_Wire_0[72]);
  not KeyNOTGate_0_37(N1815, KeyNOTWire_0[37]);
  nor NOR2_467 (keyinput_Wire_0[73], N1714, N1759);
  xor keyGate_0_73(N1819, keyinput73, keyinput_Wire_0[73]);
  nor NOR2_468 (keyinput_Wire_0[74], N1759, N1221);
  xor keyGate_0_74(KeyNOTWire_0[38], keyinput74, keyinput_Wire_0[74]);
  not KeyNOTGate_0_38(N1820, KeyNOTWire_0[38]);
  nor NOR2_469 (keyinput_Wire_0[75], N1624, N1759);
  xor keyGate_0_75(N1821, keyinput75, keyinput_Wire_0[75]);
nor NOR2_470 (N1824, N1717, N1763);
nor NOR2_471 (N1825, N1763, N549);
nor NOR2_472 (N1826, N1628, N1763);
nor NOR2_473 (N1829, N1720, N1767);
nor NOR2_474 (N1830, N1767, N597);
nor NOR2_475 (N1831, N1632, N1767);
nor NOR2_476 (N1834, N1723, N1771);
nor NOR2_477 (N1835, N1771, N645);
nor NOR2_478 (N1836, N1636, N1771);
nor NOR2_479 (N1839, N1726, N1775);
nor NOR2_480 (N1840, N1775, N693);
nor NOR2_481 (N1841, N1640, N1775);
nor NOR2_482 (N1844, N1729, N1779);
nor NOR2_483 (N1845, N1779, N741);
nor NOR2_484 (N1846, N1644, N1779);
nor NOR2_485 (N1849, N1732, N1783);
nor NOR2_486 (N1850, N1783, N789);
nor NOR2_487 (N1851, N1648, N1783);
nor NOR2_488 (N1854, N1735, N1787);
nor NOR2_489 (N1855, N1787, N837);
nor NOR2_490 (N1856, N1652, N1787);
nor NOR2_491 (N1859, N1738, N1791);
nor NOR2_492 (N1860, N1791, N885);
nor NOR2_493 (N1861, N1656, N1791);
nor NOR2_494 (N1864, N1741, N1795);
nor NOR2_495 (N1865, N1795, N933);
nor NOR2_496 (N1866, N1660, N1795);
nor NOR2_497 (N1869, N1744, N1799);
nor NOR2_498 (N1870, N1799, N981);
nor NOR2_499 (N1871, N1664, N1799);
nor NOR2_500 (N1874, N1747, N1803);
nor NOR2_501 (N1875, N1803, N1029);
nor NOR2_502 (N1876, N1668, N1803);
nor NOR2_503 (N1879, N1750, N1807);
nor NOR2_504 (N1880, N1807, N1077);
nor NOR2_505 (N1881, N1672, N1807);
nor NOR2_506 (N1884, N1753, N1811);
nor NOR2_507 (N1885, N1811, N1125);
nor NOR2_508 (N1886, N1676, N1811);
nor NOR2_509 (N1889, N1756, N1815);
nor NOR2_510 (N1890, N1815, N1173);
  nor NOR2_511 (keyinput_Wire_0[76], N1680, N1815);
  xnor keyGate_0_76(N1891, keyinput76, keyinput_Wire_0[76]);
  nor NOR2_512 (keyinput_Wire_0[77], N1819, N1820);
  xnor keyGate_0_77(KeyNOTWire_0[39], keyinput77, keyinput_Wire_0[77]);
  not KeyNOTGate_0_39(N1894, KeyNOTWire_0[39]);
  nor NOR2_513 (keyinput_Wire_0[78], N1269, N1821);
  xor keyGate_0_78(N1897, keyinput78, keyinput_Wire_0[78]);
nor NOR2_514 (N1901, N1824, N1825);
nor NOR2_515 (N1902, N1829, N1830);
nor NOR2_516 (N1905, N1834, N1835);
nor NOR2_517 (N1908, N1839, N1840);
nor NOR2_518 (N1911, N1844, N1845);
nor NOR2_519 (N1914, N1849, N1850);
nor NOR2_520 (N1917, N1854, N1855);
nor NOR2_521 (N1920, N1859, N1860);
nor NOR2_522 (N1923, N1864, N1865);
nor NOR2_523 (N1926, N1869, N1870);
nor NOR2_524 (N1929, N1874, N1875);
nor NOR2_525 (N1932, N1879, N1880);
nor NOR2_526 (N1935, N1884, N1885);
nor NOR2_527 (N1938, N1889, N1890);
  nor NOR2_528 (keyinput_Wire_0[79], N1894, N1891);
  xnor keyGate_0_79(KeyNOTWire_0[40], keyinput79, keyinput_Wire_0[79]);
  not KeyNOTGate_0_40(N1941, KeyNOTWire_0[40]);
  nor NOR2_529 (keyinput_Wire_0[80], N1269, N1897);
  xor keyGate_0_80(N1945, keyinput80, keyinput_Wire_0[80]);
  nor NOR2_530 (keyinput_Wire_0[81], N1897, N1821);
  xnor keyGate_0_81(KeyNOTWire_0[41], keyinput81, keyinput_Wire_0[81]);
  not KeyNOTGate_0_41(N1946, KeyNOTWire_0[41]);
nor NOR2_531 (N1947, N1902, N1826);
nor NOR2_532 (N1951, N1905, N1831);
nor NOR2_533 (N1955, N1908, N1836);
nor NOR2_534 (N1959, N1911, N1841);
nor NOR2_535 (N1963, N1914, N1846);
nor NOR2_536 (N1967, N1917, N1851);
nor NOR2_537 (N1971, N1920, N1856);
nor NOR2_538 (N1975, N1923, N1861);
nor NOR2_539 (N1979, N1926, N1866);
nor NOR2_540 (N1983, N1929, N1871);
nor NOR2_541 (N1987, N1932, N1876);
nor NOR2_542 (N1991, N1935, N1881);
nor NOR2_543 (N1995, N1938, N1886);
  nor NOR2_544 (keyinput_Wire_0[82], N1894, N1941);
  xor keyGate_0_82(KeyNOTWire_0[42], keyinput82, keyinput_Wire_0[82]);
  not KeyNOTGate_0_42(N1999, KeyNOTWire_0[42]);
  nor NOR2_545 (keyinput_Wire_0[83], N1941, N1891);
  xor keyGate_0_83(KeyNOTWire_0[43], keyinput83, keyinput_Wire_0[83]);
  not KeyNOTGate_0_43(N2000, KeyNOTWire_0[43]);
  nor NOR2_546 (keyinput_Wire_0[84], N1945, N1946);
  xnor keyGate_0_84(KeyNOTWire_0[44], keyinput84, keyinput_Wire_0[84]);
  not KeyNOTGate_0_44(N2001, KeyNOTWire_0[44]);
nor NOR2_547 (N2004, N1902, N1947);
nor NOR2_548 (N2005, N1947, N1826);
nor NOR2_549 (N2006, N1905, N1951);
nor NOR2_550 (N2007, N1951, N1831);
nor NOR2_551 (N2008, N1908, N1955);
nor NOR2_552 (N2009, N1955, N1836);
nor NOR2_553 (N2010, N1911, N1959);
nor NOR2_554 (N2011, N1959, N1841);
nor NOR2_555 (N2012, N1914, N1963);
nor NOR2_556 (N2013, N1963, N1846);
nor NOR2_557 (N2014, N1917, N1967);
nor NOR2_558 (N2015, N1967, N1851);
nor NOR2_559 (N2016, N1920, N1971);
nor NOR2_560 (N2017, N1971, N1856);
nor NOR2_561 (N2018, N1923, N1975);
nor NOR2_562 (N2019, N1975, N1861);
nor NOR2_563 (N2020, N1926, N1979);
nor NOR2_564 (N2021, N1979, N1866);
nor NOR2_565 (N2022, N1929, N1983);
nor NOR2_566 (N2023, N1983, N1871);
nor NOR2_567 (N2024, N1932, N1987);
nor NOR2_568 (N2025, N1987, N1876);
nor NOR2_569 (N2026, N1935, N1991);
nor NOR2_570 (N2027, N1991, N1881);
nor NOR2_571 (N2028, N1938, N1995);
nor NOR2_572 (N2029, N1995, N1886);
  nor NOR2_573 (keyinput_Wire_0[85], N1999, N2000);
  xor keyGate_0_85(KeyNOTWire_0[45], keyinput85, keyinput_Wire_0[85]);
  not KeyNOTGate_0_45(N2030, KeyNOTWire_0[45]);
  nor NOR2_574 (keyinput_Wire_0[86], N2001, N1224);
  xnor keyGate_0_86(N2033, keyinput86, keyinput_Wire_0[86]);
nor NOR2_575 (N2037, N2004, N2005);
nor NOR2_576 (N2040, N2006, N2007);
nor NOR2_577 (N2043, N2008, N2009);
nor NOR2_578 (N2046, N2010, N2011);
nor NOR2_579 (N2049, N2012, N2013);
nor NOR2_580 (N2052, N2014, N2015);
nor NOR2_581 (N2055, N2016, N2017);
nor NOR2_582 (N2058, N2018, N2019);
nor NOR2_583 (N2061, N2020, N2021);
nor NOR2_584 (N2064, N2022, N2023);
nor NOR2_585 (N2067, N2024, N2025);
nor NOR2_586 (N2070, N2026, N2027);
nor NOR2_587 (N2073, N2028, N2029);
  nor NOR2_588 (keyinput_Wire_0[87], N2030, N1176);
  xor keyGate_0_87(KeyNOTWire_0[46], keyinput87, keyinput_Wire_0[87]);
  not KeyNOTGate_0_46(N2076, KeyNOTWire_0[46]);
  nor NOR2_589 (keyinput_Wire_0[88], N2001, N2033);
  xor keyGate_0_88(KeyNOTWire_0[47], keyinput88, keyinput_Wire_0[88]);
  not KeyNOTGate_0_47(N2080, KeyNOTWire_0[47]);
  nor NOR2_590 (keyinput_Wire_0[89], N2033, N1224);
  xor keyGate_0_89(KeyNOTWire_0[48], keyinput89, keyinput_Wire_0[89]);
  not KeyNOTGate_0_48(N2081, KeyNOTWire_0[48]);
  nor NOR2_591 (keyinput_Wire_0[90], N1897, N2033);
  xnor keyGate_0_90(N2082, keyinput90, keyinput_Wire_0[90]);
nor NOR2_592 (N2085, N2037, N552);
nor NOR2_593 (N2089, N2040, N600);
nor NOR2_594 (N2093, N2043, N648);
nor NOR2_595 (N2097, N2046, N696);
nor NOR2_596 (N2101, N2049, N744);
nor NOR2_597 (N2105, N2052, N792);
nor NOR2_598 (N2109, N2055, N840);
nor NOR2_599 (N2113, N2058, N888);
nor NOR2_600 (N2117, N2061, N936);
nor NOR2_601 (N2121, N2064, N984);
nor NOR2_602 (N2125, N2067, N1032);
nor NOR2_603 (N2129, N2070, N1080);
nor NOR2_604 (N2133, N2073, N1128);
nor NOR2_605 (N2137, N2030, N2076);
nor NOR2_606 (N2138, N2076, N1176);
  nor NOR2_607 (keyinput_Wire_0[91], N1941, N2076);
  xnor keyGate_0_91(KeyNOTWire_0[49], keyinput91, keyinput_Wire_0[91]);
  not KeyNOTGate_0_49(N2139, KeyNOTWire_0[49]);
  nor NOR2_608 (keyinput_Wire_0[92], N2080, N2081);
  xnor keyGate_0_92(KeyNOTWire_0[50], keyinput92, keyinput_Wire_0[92]);
  not KeyNOTGate_0_50(N2142, KeyNOTWire_0[50]);
  nor NOR2_609 (keyinput_Wire_0[93], N1272, N2082);
  xor keyGate_0_93(KeyNOTWire_0[51], keyinput93, keyinput_Wire_0[93]);
  not KeyNOTGate_0_51(N2145, KeyNOTWire_0[51]);
nor NOR2_610 (N2149, N2037, N2085);
nor NOR2_611 (N2150, N2085, N552);
nor NOR2_612 (N2151, N1947, N2085);
nor NOR2_613 (N2154, N2040, N2089);
nor NOR2_614 (N2155, N2089, N600);
nor NOR2_615 (N2156, N1951, N2089);
nor NOR2_616 (N2159, N2043, N2093);
nor NOR2_617 (N2160, N2093, N648);
nor NOR2_618 (N2161, N1955, N2093);
nor NOR2_619 (N2164, N2046, N2097);
nor NOR2_620 (N2165, N2097, N696);
nor NOR2_621 (N2166, N1959, N2097);
nor NOR2_622 (N2169, N2049, N2101);
nor NOR2_623 (N2170, N2101, N744);
nor NOR2_624 (N2171, N1963, N2101);
nor NOR2_625 (N2174, N2052, N2105);
nor NOR2_626 (N2175, N2105, N792);
nor NOR2_627 (N2176, N1967, N2105);
nor NOR2_628 (N2179, N2055, N2109);
nor NOR2_629 (N2180, N2109, N840);
nor NOR2_630 (N2181, N1971, N2109);
nor NOR2_631 (N2184, N2058, N2113);
nor NOR2_632 (N2185, N2113, N888);
nor NOR2_633 (N2186, N1975, N2113);
nor NOR2_634 (N2189, N2061, N2117);
nor NOR2_635 (N2190, N2117, N936);
nor NOR2_636 (N2191, N1979, N2117);
nor NOR2_637 (N2194, N2064, N2121);
nor NOR2_638 (N2195, N2121, N984);
nor NOR2_639 (N2196, N1983, N2121);
nor NOR2_640 (N2199, N2067, N2125);
nor NOR2_641 (N2200, N2125, N1032);
nor NOR2_642 (N2201, N1987, N2125);
nor NOR2_643 (N2204, N2070, N2129);
nor NOR2_644 (N2205, N2129, N1080);
nor NOR2_645 (N2206, N1991, N2129);
nor NOR2_646 (N2209, N2073, N2133);
nor NOR2_647 (N2210, N2133, N1128);
nor NOR2_648 (N2211, N1995, N2133);
nor NOR2_649 (N2214, N2137, N2138);
  nor NOR2_650 (keyinput_Wire_0[94], N2142, N2139);
  xor keyGate_0_94(N2217, keyinput94, keyinput_Wire_0[94]);
  nor NOR2_651 (keyinput_Wire_0[95], N1272, N2145);
  xnor keyGate_0_95(KeyNOTWire_0[52], keyinput95, keyinput_Wire_0[95]);
  not KeyNOTGate_0_52(N2221, KeyNOTWire_0[52]);
  nor NOR2_652 (keyinput_Wire_0[96], N2145, N2082);
  xor keyGate_0_96(N2222, keyinput96, keyinput_Wire_0[96]);
nor NOR2_653 (N2223, N2149, N2150);
nor NOR2_654 (N2224, N2154, N2155);
nor NOR2_655 (N2227, N2159, N2160);
nor NOR2_656 (N2230, N2164, N2165);
nor NOR2_657 (N2233, N2169, N2170);
nor NOR2_658 (N2236, N2174, N2175);
nor NOR2_659 (N2239, N2179, N2180);
nor NOR2_660 (N2242, N2184, N2185);
nor NOR2_661 (N2245, N2189, N2190);
nor NOR2_662 (N2248, N2194, N2195);
nor NOR2_663 (N2251, N2199, N2200);
nor NOR2_664 (N2254, N2204, N2205);
nor NOR2_665 (N2257, N2209, N2210);
nor NOR2_666 (N2260, N2214, N2211);
  nor NOR2_667 (keyinput_Wire_0[97], N2142, N2217);
  xnor keyGate_0_97(KeyNOTWire_0[53], keyinput97, keyinput_Wire_0[97]);
  not KeyNOTGate_0_53(N2264, KeyNOTWire_0[53]);
  nor NOR2_668 (keyinput_Wire_0[98], N2217, N2139);
  xnor keyGate_0_98(KeyNOTWire_0[54], keyinput98, keyinput_Wire_0[98]);
  not KeyNOTGate_0_54(N2265, KeyNOTWire_0[54]);
  nor NOR2_669 (keyinput_Wire_0[99], N2221, N2222);
  xnor keyGate_0_99(N2266, keyinput99, keyinput_Wire_0[99]);
nor NOR2_670 (N2269, N2224, N2151);
nor NOR2_671 (N2273, N2227, N2156);
nor NOR2_672 (N2277, N2230, N2161);
nor NOR2_673 (N2281, N2233, N2166);
nor NOR2_674 (N2285, N2236, N2171);
nor NOR2_675 (N2289, N2239, N2176);
nor NOR2_676 (N2293, N2242, N2181);
nor NOR2_677 (N2297, N2245, N2186);
nor NOR2_678 (N2301, N2248, N2191);
nor NOR2_679 (N2305, N2251, N2196);
nor NOR2_680 (N2309, N2254, N2201);
nor NOR2_681 (N2313, N2257, N2206);
nor NOR2_682 (N2317, N2214, N2260);
nor NOR2_683 (N2318, N2260, N2211);
  nor NOR2_684 (keyinput_Wire_0[100], N2264, N2265);
  xor keyGate_0_100(N2319, keyinput100, keyinput_Wire_0[100]);
  nor NOR2_685 (keyinput_Wire_0[101], N2266, N1227);
  xor keyGate_0_101(KeyNOTWire_0[55], keyinput101, keyinput_Wire_0[101]);
  not KeyNOTGate_0_55(N2322, KeyNOTWire_0[55]);
nor NOR2_686 (N2326, N2224, N2269);
nor NOR2_687 (N2327, N2269, N2151);
nor NOR2_688 (N2328, N2227, N2273);
nor NOR2_689 (N2329, N2273, N2156);
nor NOR2_690 (N2330, N2230, N2277);
nor NOR2_691 (N2331, N2277, N2161);
  nor NOR2_692 (keyinput_Wire_0[102], N2233, N2281);
  xor keyGate_0_102(KeyNOTWire_0[56], keyinput102, keyinput_Wire_0[102]);
  not KeyNOTGate_0_56(N2332, KeyNOTWire_0[56]);
nor NOR2_693 (N2333, N2281, N2166);
nor NOR2_694 (N2334, N2236, N2285);
nor NOR2_695 (N2335, N2285, N2171);
nor NOR2_696 (N2336, N2239, N2289);
nor NOR2_697 (N2337, N2289, N2176);
nor NOR2_698 (N2338, N2242, N2293);
nor NOR2_699 (N2339, N2293, N2181);
nor NOR2_700 (N2340, N2245, N2297);
nor NOR2_701 (N2341, N2297, N2186);
nor NOR2_702 (N2342, N2248, N2301);
nor NOR2_703 (N2343, N2301, N2191);
nor NOR2_704 (N2344, N2251, N2305);
nor NOR2_705 (N2345, N2305, N2196);
nor NOR2_706 (N2346, N2254, N2309);
nor NOR2_707 (N2347, N2309, N2201);
nor NOR2_708 (N2348, N2257, N2313);
nor NOR2_709 (N2349, N2313, N2206);
nor NOR2_710 (N2350, N2317, N2318);
  nor NOR2_711 (keyinput_Wire_0[103], N2319, N1179);
  xnor keyGate_0_103(N2353, keyinput103, keyinput_Wire_0[103]);
  nor NOR2_712 (keyinput_Wire_0[104], N2266, N2322);
  xor keyGate_0_104(KeyNOTWire_0[57], keyinput104, keyinput_Wire_0[104]);
  not KeyNOTGate_0_57(N2357, KeyNOTWire_0[57]);
  nor NOR2_713 (keyinput_Wire_0[105], N2322, N1227);
  xor keyGate_0_105(N2358, keyinput105, keyinput_Wire_0[105]);
  nor NOR2_714 (keyinput_Wire_0[106], N2145, N2322);
  xor keyGate_0_106(N2359, keyinput106, keyinput_Wire_0[106]);
nor NOR2_715 (N2362, N2326, N2327);
nor NOR2_716 (N2365, N2328, N2329);
nor NOR2_717 (N2368, N2330, N2331);
nor NOR2_718 (N2371, N2332, N2333);
nor NOR2_719 (N2374, N2334, N2335);
nor NOR2_720 (N2377, N2336, N2337);
nor NOR2_721 (N2380, N2338, N2339);
nor NOR2_722 (N2383, N2340, N2341);
nor NOR2_723 (N2386, N2342, N2343);
nor NOR2_724 (N2389, N2344, N2345);
nor NOR2_725 (N2392, N2346, N2347);
nor NOR2_726 (N2395, N2348, N2349);
nor NOR2_727 (N2398, N2350, N1131);
nor NOR2_728 (N2402, N2319, N2353);
nor NOR2_729 (N2403, N2353, N1179);
  nor NOR2_730 (keyinput_Wire_0[107], N2217, N2353);
  xnor keyGate_0_107(KeyNOTWire_0[58], keyinput107, keyinput_Wire_0[107]);
  not KeyNOTGate_0_58(N2404, KeyNOTWire_0[58]);
  nor NOR2_731 (keyinput_Wire_0[108], N2357, N2358);
  xnor keyGate_0_108(N2407, keyinput108, keyinput_Wire_0[108]);
  nor NOR2_732 (keyinput_Wire_0[109], N1275, N2359);
  xor keyGate_0_109(KeyNOTWire_0[59], keyinput109, keyinput_Wire_0[109]);
  not KeyNOTGate_0_59(N2410, KeyNOTWire_0[59]);
nor NOR2_733 (N2414, N2362, N555);
nor NOR2_734 (N2418, N2365, N603);
nor NOR2_735 (N2422, N2368, N651);
nor NOR2_736 (N2426, N2371, N699);
nor NOR2_737 (N2430, N2374, N747);
nor NOR2_738 (N2434, N2377, N795);
nor NOR2_739 (N2438, N2380, N843);
nor NOR2_740 (N2442, N2383, N891);
nor NOR2_741 (N2446, N2386, N939);
nor NOR2_742 (N2450, N2389, N987);
nor NOR2_743 (N2454, N2392, N1035);
nor NOR2_744 (N2458, N2395, N1083);
nor NOR2_745 (N2462, N2350, N2398);
nor NOR2_746 (N2463, N2398, N1131);
nor NOR2_747 (N2464, N2260, N2398);
nor NOR2_748 (N2467, N2402, N2403);
  nor NOR2_749 (keyinput_Wire_0[110], N2407, N2404);
  xor keyGate_0_110(N2470, keyinput110, keyinput_Wire_0[110]);
  nor NOR2_750 (keyinput_Wire_0[111], N1275, N2410);
  xnor keyGate_0_111(KeyNOTWire_0[60], keyinput111, keyinput_Wire_0[111]);
  not KeyNOTGate_0_60(N2474, KeyNOTWire_0[60]);
  nor NOR2_751 (keyinput_Wire_0[112], N2410, N2359);
  xor keyGate_0_112(KeyNOTWire_0[61], keyinput112, keyinput_Wire_0[112]);
  not KeyNOTGate_0_61(N2475, KeyNOTWire_0[61]);
nor NOR2_752 (N2476, N2362, N2414);
nor NOR2_753 (N2477, N2414, N555);
nor NOR2_754 (N2478, N2269, N2414);
nor NOR2_755 (N2481, N2365, N2418);
nor NOR2_756 (N2482, N2418, N603);
nor NOR2_757 (N2483, N2273, N2418);
nor NOR2_758 (N2486, N2368, N2422);
nor NOR2_759 (N2487, N2422, N651);
nor NOR2_760 (N2488, N2277, N2422);
nor NOR2_761 (N2491, N2371, N2426);
nor NOR2_762 (N2492, N2426, N699);
nor NOR2_763 (N2493, N2281, N2426);
nor NOR2_764 (N2496, N2374, N2430);
nor NOR2_765 (N2497, N2430, N747);
nor NOR2_766 (N2498, N2285, N2430);
nor NOR2_767 (N2501, N2377, N2434);
nor NOR2_768 (N2502, N2434, N795);
nor NOR2_769 (N2503, N2289, N2434);
nor NOR2_770 (N2506, N2380, N2438);
nor NOR2_771 (N2507, N2438, N843);
nor NOR2_772 (N2508, N2293, N2438);
nor NOR2_773 (N2511, N2383, N2442);
nor NOR2_774 (N2512, N2442, N891);
nor NOR2_775 (N2513, N2297, N2442);
nor NOR2_776 (N2516, N2386, N2446);
nor NOR2_777 (N2517, N2446, N939);
nor NOR2_778 (N2518, N2301, N2446);
nor NOR2_779 (N2521, N2389, N2450);
nor NOR2_780 (N2522, N2450, N987);
nor NOR2_781 (N2523, N2305, N2450);
nor NOR2_782 (N2526, N2392, N2454);
nor NOR2_783 (N2527, N2454, N1035);
nor NOR2_784 (N2528, N2309, N2454);
nor NOR2_785 (N2531, N2395, N2458);
nor NOR2_786 (N2532, N2458, N1083);
nor NOR2_787 (N2533, N2313, N2458);
nor NOR2_788 (N2536, N2462, N2463);
nor NOR2_789 (N2539, N2467, N2464);
  nor NOR2_790 (keyinput_Wire_0[113], N2407, N2470);
  xor keyGate_0_113(KeyNOTWire_0[62], keyinput113, keyinput_Wire_0[113]);
  not KeyNOTGate_0_62(N2543, KeyNOTWire_0[62]);
  nor NOR2_791 (keyinput_Wire_0[114], N2470, N2404);
  xor keyGate_0_114(KeyNOTWire_0[63], keyinput114, keyinput_Wire_0[114]);
  not KeyNOTGate_0_63(N2544, KeyNOTWire_0[63]);
  nor NOR2_792 (keyinput_Wire_0[115], N2474, N2475);
  xor keyGate_0_115(N2545, keyinput115, keyinput_Wire_0[115]);
nor NOR2_793 (N2548, N2476, N2477);
nor NOR2_794 (N2549, N2481, N2482);
nor NOR2_795 (N2552, N2486, N2487);
nor NOR2_796 (N2555, N2491, N2492);
nor NOR2_797 (N2558, N2496, N2497);
nor NOR2_798 (N2561, N2501, N2502);
nor NOR2_799 (N2564, N2506, N2507);
nor NOR2_800 (N2567, N2511, N2512);
nor NOR2_801 (N2570, N2516, N2517);
nor NOR2_802 (N2573, N2521, N2522);
nor NOR2_803 (N2576, N2526, N2527);
nor NOR2_804 (N2579, N2531, N2532);
nor NOR2_805 (N2582, N2536, N2533);
nor NOR2_806 (N2586, N2467, N2539);
nor NOR2_807 (N2587, N2539, N2464);
  nor NOR2_808 (keyinput_Wire_0[116], N2543, N2544);
  xor keyGate_0_116(N2588, keyinput116, keyinput_Wire_0[116]);
  nor NOR2_809 (keyinput_Wire_0[117], N2545, N1230);
  xor keyGate_0_117(KeyNOTWire_0[64], keyinput117, keyinput_Wire_0[117]);
  not KeyNOTGate_0_64(N2591, KeyNOTWire_0[64]);
nor NOR2_810 (N2595, N2549, N2478);
nor NOR2_811 (N2599, N2552, N2483);
nor NOR2_812 (N2603, N2555, N2488);
  nor NOR2_813 (keyinput_Wire_0[118], N2558, N2493);
  xnor keyGate_0_118(KeyNOTWire_0[65], keyinput118, keyinput_Wire_0[118]);
  not KeyNOTGate_0_65(N2607, KeyNOTWire_0[65]);
nor NOR2_814 (N2611, N2561, N2498);
nor NOR2_815 (N2615, N2564, N2503);
nor NOR2_816 (N2619, N2567, N2508);
nor NOR2_817 (N2623, N2570, N2513);
nor NOR2_818 (N2627, N2573, N2518);
nor NOR2_819 (N2631, N2576, N2523);
nor NOR2_820 (N2635, N2579, N2528);
nor NOR2_821 (N2639, N2536, N2582);
nor NOR2_822 (N2640, N2582, N2533);
nor NOR2_823 (N2641, N2586, N2587);
  nor NOR2_824 (keyinput_Wire_0[119], N2588, N1182);
  xnor keyGate_0_119(KeyNOTWire_0[66], keyinput119, keyinput_Wire_0[119]);
  not KeyNOTGate_0_66(N2644, KeyNOTWire_0[66]);
  nor NOR2_825 (keyinput_Wire_0[120], N2545, N2591);
  xnor keyGate_0_120(KeyNOTWire_0[67], keyinput120, keyinput_Wire_0[120]);
  not KeyNOTGate_0_67(N2648, KeyNOTWire_0[67]);
  nor NOR2_826 (keyinput_Wire_0[121], N2591, N1230);
  xnor keyGate_0_121(N2649, keyinput121, keyinput_Wire_0[121]);
  nor NOR2_827 (keyinput_Wire_0[122], N2410, N2591);
  xnor keyGate_0_122(KeyNOTWire_0[68], keyinput122, keyinput_Wire_0[122]);
  not KeyNOTGate_0_68(N2650, KeyNOTWire_0[68]);
nor NOR2_828 (N2653, N2549, N2595);
nor NOR2_829 (N2654, N2595, N2478);
nor NOR2_830 (N2655, N2552, N2599);
nor NOR2_831 (N2656, N2599, N2483);
nor NOR2_832 (N2657, N2555, N2603);
nor NOR2_833 (N2658, N2603, N2488);
nor NOR2_834 (N2659, N2558, N2607);
nor NOR2_835 (N2660, N2607, N2493);
nor NOR2_836 (N2661, N2561, N2611);
nor NOR2_837 (N2662, N2611, N2498);
nor NOR2_838 (N2663, N2564, N2615);
nor NOR2_839 (N2664, N2615, N2503);
nor NOR2_840 (N2665, N2567, N2619);
nor NOR2_841 (N2666, N2619, N2508);
nor NOR2_842 (N2667, N2570, N2623);
nor NOR2_843 (N2668, N2623, N2513);
nor NOR2_844 (N2669, N2573, N2627);
nor NOR2_845 (N2670, N2627, N2518);
nor NOR2_846 (N2671, N2576, N2631);
nor NOR2_847 (N2672, N2631, N2523);
nor NOR2_848 (N2673, N2579, N2635);
nor NOR2_849 (N2674, N2635, N2528);
nor NOR2_850 (N2675, N2639, N2640);
nor NOR2_851 (N2678, N2641, N1134);
nor NOR2_852 (N2682, N2588, N2644);
nor NOR2_853 (N2683, N2644, N1182);
  nor NOR2_854 (keyinput_Wire_0[123], N2470, N2644);
  xnor keyGate_0_123(KeyNOTWire_0[69], keyinput123, keyinput_Wire_0[123]);
  not KeyNOTGate_0_69(N2684, KeyNOTWire_0[69]);
  nor NOR2_855 (keyinput_Wire_0[124], N2648, N2649);
  xor keyGate_0_124(KeyNOTWire_0[70], keyinput124, keyinput_Wire_0[124]);
  not KeyNOTGate_0_70(N2687, KeyNOTWire_0[70]);
  nor NOR2_856 (keyinput_Wire_0[125], N1278, N2650);
  xor keyGate_0_125(N2690, keyinput125, keyinput_Wire_0[125]);
nor NOR2_857 (N2694, N2653, N2654);
nor NOR2_858 (N2697, N2655, N2656);
nor NOR2_859 (N2700, N2657, N2658);
nor NOR2_860 (N2703, N2659, N2660);
nor NOR2_861 (N2706, N2661, N2662);
nor NOR2_862 (N2709, N2663, N2664);
nor NOR2_863 (N2712, N2665, N2666);
nor NOR2_864 (N2715, N2667, N2668);
nor NOR2_865 (N2718, N2669, N2670);
nor NOR2_866 (N2721, N2671, N2672);
nor NOR2_867 (N2724, N2673, N2674);
nor NOR2_868 (N2727, N2675, N1086);
nor NOR2_869 (N2731, N2641, N2678);
nor NOR2_870 (N2732, N2678, N1134);
nor NOR2_871 (N2733, N2539, N2678);
nor NOR2_872 (N2736, N2682, N2683);
  nor NOR2_873 (keyinput_Wire_0[126], N2687, N2684);
  xor keyGate_0_126(N2739, keyinput126, keyinput_Wire_0[126]);
  nor NOR2_874 (keyinput_Wire_0[127], N1278, N2690);
  xor keyGate_0_127(KeyNOTWire_0[71], keyinput127, keyinput_Wire_0[127]);
  not KeyNOTGate_0_71(N2743, KeyNOTWire_0[71]);
  nor NOR2_875 (keyinput_Wire_0[128], N2690, N2650);
  xnor keyGate_0_128(KeyNOTWire_0[72], keyinput128, keyinput_Wire_0[128]);
  not KeyNOTGate_0_72(N2744, KeyNOTWire_0[72]);
nor NOR2_876 (N2745, N2694, N558);
nor NOR2_877 (N2749, N2697, N606);
nor NOR2_878 (N2753, N2700, N654);
nor NOR2_879 (N2757, N2703, N702);
nor NOR2_880 (N2761, N2706, N750);
nor NOR2_881 (N2765, N2709, N798);
nor NOR2_882 (N2769, N2712, N846);
nor NOR2_883 (N2773, N2715, N894);
nor NOR2_884 (N2777, N2718, N942);
nor NOR2_885 (N2781, N2721, N990);
nor NOR2_886 (N2785, N2724, N1038);
nor NOR2_887 (N2789, N2675, N2727);
nor NOR2_888 (N2790, N2727, N1086);
nor NOR2_889 (N2791, N2582, N2727);
nor NOR2_890 (N2794, N2731, N2732);
nor NOR2_891 (N2797, N2736, N2733);
  nor NOR2_892 (keyinput_Wire_0[129], N2687, N2739);
  xor keyGate_0_129(N2801, keyinput129, keyinput_Wire_0[129]);
  nor NOR2_893 (keyinput_Wire_0[130], N2739, N2684);
  xor keyGate_0_130(N2802, keyinput130, keyinput_Wire_0[130]);
  nor NOR2_894 (keyinput_Wire_0[131], N2743, N2744);
  xnor keyGate_0_131(N2803, keyinput131, keyinput_Wire_0[131]);
nor NOR2_895 (N2806, N2694, N2745);
nor NOR2_896 (N2807, N2745, N558);
nor NOR2_897 (N2808, N2595, N2745);
nor NOR2_898 (N2811, N2697, N2749);
nor NOR2_899 (N2812, N2749, N606);
nor NOR2_900 (N2813, N2599, N2749);
nor NOR2_901 (N2816, N2700, N2753);
nor NOR2_902 (N2817, N2753, N654);
nor NOR2_903 (N2818, N2603, N2753);
nor NOR2_904 (N2821, N2703, N2757);
nor NOR2_905 (N2822, N2757, N702);
nor NOR2_906 (N2823, N2607, N2757);
nor NOR2_907 (N2826, N2706, N2761);
nor NOR2_908 (N2827, N2761, N750);
nor NOR2_909 (N2828, N2611, N2761);
nor NOR2_910 (N2831, N2709, N2765);
nor NOR2_911 (N2832, N2765, N798);
nor NOR2_912 (N2833, N2615, N2765);
nor NOR2_913 (N2836, N2712, N2769);
nor NOR2_914 (N2837, N2769, N846);
nor NOR2_915 (N2838, N2619, N2769);
nor NOR2_916 (N2841, N2715, N2773);
nor NOR2_917 (N2842, N2773, N894);
nor NOR2_918 (N2843, N2623, N2773);
nor NOR2_919 (N2846, N2718, N2777);
nor NOR2_920 (N2847, N2777, N942);
nor NOR2_921 (N2848, N2627, N2777);
nor NOR2_922 (N2851, N2721, N2781);
nor NOR2_923 (N2852, N2781, N990);
nor NOR2_924 (N2853, N2631, N2781);
nor NOR2_925 (N2856, N2724, N2785);
nor NOR2_926 (N2857, N2785, N1038);
nor NOR2_927 (N2858, N2635, N2785);
nor NOR2_928 (N2861, N2789, N2790);
nor NOR2_929 (N2864, N2794, N2791);
nor NOR2_930 (N2868, N2736, N2797);
nor NOR2_931 (N2869, N2797, N2733);
  nor NOR2_932 (keyinput_Wire_0[132], N2801, N2802);
  xnor keyGate_0_132(N2870, keyinput132, keyinput_Wire_0[132]);
  nor NOR2_933 (keyinput_Wire_0[133], N2803, N1233);
  xnor keyGate_0_133(N2873, keyinput133, keyinput_Wire_0[133]);
nor NOR2_934 (N2877, N2806, N2807);
nor NOR2_935 (N2878, N2811, N2812);
nor NOR2_936 (N2881, N2816, N2817);
nor NOR2_937 (N2884, N2821, N2822);
nor NOR2_938 (N2887, N2826, N2827);
nor NOR2_939 (N2890, N2831, N2832);
nor NOR2_940 (N2893, N2836, N2837);
nor NOR2_941 (N2896, N2841, N2842);
nor NOR2_942 (N2899, N2846, N2847);
nor NOR2_943 (N2902, N2851, N2852);
nor NOR2_944 (N2905, N2856, N2857);
nor NOR2_945 (N2908, N2861, N2858);
nor NOR2_946 (N2912, N2794, N2864);
nor NOR2_947 (N2913, N2864, N2791);
nor NOR2_948 (N2914, N2868, N2869);
  nor NOR2_949 (keyinput_Wire_0[134], N2870, N1185);
  xor keyGate_0_134(KeyNOTWire_0[73], keyinput134, keyinput_Wire_0[134]);
  not KeyNOTGate_0_73(N2917, KeyNOTWire_0[73]);
  nor NOR2_950 (keyinput_Wire_0[135], N2803, N2873);
  xor keyGate_0_135(N2921, keyinput135, keyinput_Wire_0[135]);
  nor NOR2_951 (keyinput_Wire_0[136], N2873, N1233);
  xor keyGate_0_136(KeyNOTWire_0[74], keyinput136, keyinput_Wire_0[136]);
  not KeyNOTGate_0_74(N2922, KeyNOTWire_0[74]);
  nor NOR2_952 (keyinput_Wire_0[137], N2690, N2873);
  xor keyGate_0_137(N2923, keyinput137, keyinput_Wire_0[137]);
nor NOR2_953 (N2926, N2878, N2808);
nor NOR2_954 (N2930, N2881, N2813);
nor NOR2_955 (N2934, N2884, N2818);
nor NOR2_956 (N2938, N2887, N2823);
nor NOR2_957 (N2942, N2890, N2828);
nor NOR2_958 (N2946, N2893, N2833);
nor NOR2_959 (N2950, N2896, N2838);
nor NOR2_960 (N2954, N2899, N2843);
nor NOR2_961 (N2958, N2902, N2848);
nor NOR2_962 (N2962, N2905, N2853);
nor NOR2_963 (N2966, N2861, N2908);
nor NOR2_964 (N2967, N2908, N2858);
nor NOR2_965 (N2968, N2912, N2913);
nor NOR2_966 (N2971, N2914, N1137);
nor NOR2_967 (N2975, N2870, N2917);
nor NOR2_968 (N2976, N2917, N1185);
  nor NOR2_969 (keyinput_Wire_0[138], N2739, N2917);
  xnor keyGate_0_138(KeyNOTWire_0[75], keyinput138, keyinput_Wire_0[138]);
  not KeyNOTGate_0_75(N2977, KeyNOTWire_0[75]);
  nor NOR2_970 (keyinput_Wire_0[139], N2921, N2922);
  xnor keyGate_0_139(N2980, keyinput139, keyinput_Wire_0[139]);
  nor NOR2_971 (keyinput_Wire_0[140], N1281, N2923);
  xor keyGate_0_140(KeyNOTWire_0[76], keyinput140, keyinput_Wire_0[140]);
  not KeyNOTGate_0_76(N2983, KeyNOTWire_0[76]);
nor NOR2_972 (N2987, N2878, N2926);
nor NOR2_973 (N2988, N2926, N2808);
nor NOR2_974 (N2989, N2881, N2930);
nor NOR2_975 (N2990, N2930, N2813);
nor NOR2_976 (N2991, N2884, N2934);
nor NOR2_977 (N2992, N2934, N2818);
nor NOR2_978 (N2993, N2887, N2938);
nor NOR2_979 (N2994, N2938, N2823);
nor NOR2_980 (N2995, N2890, N2942);
nor NOR2_981 (N2996, N2942, N2828);
nor NOR2_982 (N2997, N2893, N2946);
nor NOR2_983 (N2998, N2946, N2833);
nor NOR2_984 (N2999, N2896, N2950);
nor NOR2_985 (N3000, N2950, N2838);
nor NOR2_986 (N3001, N2899, N2954);
nor NOR2_987 (N3002, N2954, N2843);
nor NOR2_988 (N3003, N2902, N2958);
nor NOR2_989 (N3004, N2958, N2848);
nor NOR2_990 (N3005, N2905, N2962);
nor NOR2_991 (N3006, N2962, N2853);
nor NOR2_992 (N3007, N2966, N2967);
nor NOR2_993 (N3010, N2968, N1089);
nor NOR2_994 (N3014, N2914, N2971);
nor NOR2_995 (N3015, N2971, N1137);
nor NOR2_996 (N3016, N2797, N2971);
nor NOR2_997 (N3019, N2975, N2976);
  nor NOR2_998 (keyinput_Wire_0[141], N2980, N2977);
  xnor keyGate_0_141(N3022, keyinput141, keyinput_Wire_0[141]);
  nor NOR2_999 (keyinput_Wire_0[142], N1281, N2983);
  xnor keyGate_0_142(N3026, keyinput142, keyinput_Wire_0[142]);
  nor NOR2_1000 (keyinput_Wire_0[143], N2983, N2923);
  xor keyGate_0_143(N3027, keyinput143, keyinput_Wire_0[143]);
  nor NOR2_1001 (keyinput_Wire_0[144], N2987, N2988);
  xor keyGate_0_144(N3028, keyinput144, keyinput_Wire_0[144]);
nor NOR2_1002 (N3031, N2989, N2990);
nor NOR2_1003 (N3034, N2991, N2992);
nor NOR2_1004 (N3037, N2993, N2994);
nor NOR2_1005 (N3040, N2995, N2996);
nor NOR2_1006 (N3043, N2997, N2998);
nor NOR2_1007 (N3046, N2999, N3000);
nor NOR2_1008 (N3049, N3001, N3002);
nor NOR2_1009 (N3052, N3003, N3004);
nor NOR2_1010 (N3055, N3005, N3006);
nor NOR2_1011 (N3058, N3007, N1041);
nor NOR2_1012 (N3062, N2968, N3010);
nor NOR2_1013 (N3063, N3010, N1089);
nor NOR2_1014 (N3064, N2864, N3010);
nor NOR2_1015 (N3067, N3014, N3015);
nor NOR2_1016 (N3070, N3019, N3016);
  nor NOR2_1017 (keyinput_Wire_0[145], N2980, N3022);
  xor keyGate_0_145(N3074, keyinput145, keyinput_Wire_0[145]);
  nor NOR2_1018 (keyinput_Wire_0[146], N3022, N2977);
  xnor keyGate_0_146(N3075, keyinput146, keyinput_Wire_0[146]);
  nor NOR2_1019 (keyinput_Wire_0[147], N3026, N3027);
  xor keyGate_0_147(N3076, keyinput147, keyinput_Wire_0[147]);
nor NOR2_1020 (N3079, N3028, N561);
nor NOR2_1021 (N3083, N3031, N609);
nor NOR2_1022 (N3087, N3034, N657);
nor NOR2_1023 (N3091, N3037, N705);
nor NOR2_1024 (N3095, N3040, N753);
nor NOR2_1025 (N3099, N3043, N801);
nor NOR2_1026 (N3103, N3046, N849);
nor NOR2_1027 (N3107, N3049, N897);
nor NOR2_1028 (N3111, N3052, N945);
nor NOR2_1029 (N3115, N3055, N993);
nor NOR2_1030 (N3119, N3007, N3058);
nor NOR2_1031 (N3120, N3058, N1041);
nor NOR2_1032 (N3121, N2908, N3058);
nor NOR2_1033 (N3124, N3062, N3063);
nor NOR2_1034 (N3127, N3067, N3064);
nor NOR2_1035 (N3131, N3019, N3070);
nor NOR2_1036 (N3132, N3070, N3016);
  nor NOR2_1037 (keyinput_Wire_0[148], N3074, N3075);
  xor keyGate_0_148(N3133, keyinput148, keyinput_Wire_0[148]);
  nor NOR2_1038 (keyinput_Wire_0[149], N3076, N1236);
  xnor keyGate_0_149(KeyNOTWire_0[77], keyinput149, keyinput_Wire_0[149]);
  not KeyNOTGate_0_77(N3136, KeyNOTWire_0[77]);
nor NOR2_1039 (N3140, N3028, N3079);
nor NOR2_1040 (N3141, N3079, N561);
nor NOR2_1041 (N3142, N2926, N3079);
nor NOR2_1042 (N3145, N3031, N3083);
nor NOR2_1043 (N3146, N3083, N609);
nor NOR2_1044 (N3147, N2930, N3083);
nor NOR2_1045 (N3150, N3034, N3087);
nor NOR2_1046 (N3151, N3087, N657);
nor NOR2_1047 (N3152, N2934, N3087);
nor NOR2_1048 (N3155, N3037, N3091);
nor NOR2_1049 (N3156, N3091, N705);
nor NOR2_1050 (N3157, N2938, N3091);
nor NOR2_1051 (N3160, N3040, N3095);
nor NOR2_1052 (N3161, N3095, N753);
nor NOR2_1053 (N3162, N2942, N3095);
nor NOR2_1054 (N3165, N3043, N3099);
nor NOR2_1055 (N3166, N3099, N801);
nor NOR2_1056 (N3167, N2946, N3099);
nor NOR2_1057 (N3170, N3046, N3103);
nor NOR2_1058 (N3171, N3103, N849);
nor NOR2_1059 (N3172, N2950, N3103);
nor NOR2_1060 (N3175, N3049, N3107);
nor NOR2_1061 (N3176, N3107, N897);
nor NOR2_1062 (N3177, N2954, N3107);
nor NOR2_1063 (N3180, N3052, N3111);
nor NOR2_1064 (N3181, N3111, N945);
nor NOR2_1065 (N3182, N2958, N3111);
nor NOR2_1066 (N3185, N3055, N3115);
nor NOR2_1067 (N3186, N3115, N993);
nor NOR2_1068 (N3187, N2962, N3115);
nor NOR2_1069 (N3190, N3119, N3120);
nor NOR2_1070 (N3193, N3124, N3121);
nor NOR2_1071 (N3197, N3067, N3127);
nor NOR2_1072 (N3198, N3127, N3064);
nor NOR2_1073 (N3199, N3131, N3132);
  nor NOR2_1074 (keyinput_Wire_0[150], N3133, N1188);
  xnor keyGate_0_150(KeyNOTWire_0[78], keyinput150, keyinput_Wire_0[150]);
  not KeyNOTGate_0_78(N3202, KeyNOTWire_0[78]);
  nor NOR2_1075 (keyinput_Wire_0[151], N3076, N3136);
  xnor keyGate_0_151(N3206, keyinput151, keyinput_Wire_0[151]);
  nor NOR2_1076 (keyinput_Wire_0[152], N3136, N1236);
  xor keyGate_0_152(N3207, keyinput152, keyinput_Wire_0[152]);
  nor NOR2_1077 (keyinput_Wire_0[153], N2983, N3136);
  xor keyGate_0_153(N3208, keyinput153, keyinput_Wire_0[153]);
nor NOR2_1078 (N3211, N3140, N3141);
nor NOR2_1079 (N3212, N3145, N3146);
nor NOR2_1080 (N3215, N3150, N3151);
nor NOR2_1081 (N3218, N3155, N3156);
nor NOR2_1082 (N3221, N3160, N3161);
nor NOR2_1083 (N3224, N3165, N3166);
nor NOR2_1084 (N3227, N3170, N3171);
nor NOR2_1085 (N3230, N3175, N3176);
nor NOR2_1086 (N3233, N3180, N3181);
nor NOR2_1087 (N3236, N3185, N3186);
nor NOR2_1088 (N3239, N3190, N3187);
nor NOR2_1089 (N3243, N3124, N3193);
nor NOR2_1090 (N3244, N3193, N3121);
nor NOR2_1091 (N3245, N3197, N3198);
nor NOR2_1092 (N3248, N3199, N1140);
nor NOR2_1093 (N3252, N3133, N3202);
  nor NOR2_1094 (keyinput_Wire_0[154], N3202, N1188);
  xnor keyGate_0_154(N3253, keyinput154, keyinput_Wire_0[154]);
  nor NOR2_1095 (keyinput_Wire_0[155], N3022, N3202);
  xor keyGate_0_155(KeyNOTWire_0[79], keyinput155, keyinput_Wire_0[155]);
  not KeyNOTGate_0_79(N3254, KeyNOTWire_0[79]);
  nor NOR2_1096 (keyinput_Wire_0[156], N3206, N3207);
  xnor keyGate_0_156(N3257, keyinput156, keyinput_Wire_0[156]);
  nor NOR2_1097 (keyinput_Wire_0[157], N1284, N3208);
  xnor keyGate_0_157(N3260, keyinput157, keyinput_Wire_0[157]);
nor NOR2_1098 (N3264, N3212, N3142);
nor NOR2_1099 (N3268, N3215, N3147);
nor NOR2_1100 (N3272, N3218, N3152);
nor NOR2_1101 (N3276, N3221, N3157);
nor NOR2_1102 (N3280, N3224, N3162);
nor NOR2_1103 (N3284, N3227, N3167);
nor NOR2_1104 (N3288, N3230, N3172);
nor NOR2_1105 (N3292, N3233, N3177);
nor NOR2_1106 (N3296, N3236, N3182);
nor NOR2_1107 (N3300, N3190, N3239);
nor NOR2_1108 (N3301, N3239, N3187);
nor NOR2_1109 (N3302, N3243, N3244);
nor NOR2_1110 (N3305, N3245, N1092);
nor NOR2_1111 (N3309, N3199, N3248);
nor NOR2_1112 (N3310, N3248, N1140);
nor NOR2_1113 (N3311, N3070, N3248);
nor NOR2_1114 (N3314, N3252, N3253);
  nor NOR2_1115 (keyinput_Wire_0[158], N3257, N3254);
  xor keyGate_0_158(KeyNOTWire_0[80], keyinput158, keyinput_Wire_0[158]);
  not KeyNOTGate_0_80(N3317, KeyNOTWire_0[80]);
  nor NOR2_1116 (keyinput_Wire_0[159], N1284, N3260);
  xor keyGate_0_159(KeyNOTWire_0[81], keyinput159, keyinput_Wire_0[159]);
  not KeyNOTGate_0_81(N3321, KeyNOTWire_0[81]);
  nor NOR2_1117 (keyinput_Wire_0[160], N3260, N3208);
  xnor keyGate_0_160(N3322, keyinput160, keyinput_Wire_0[160]);
nor NOR2_1118 (N3323, N3212, N3264);
nor NOR2_1119 (N3324, N3264, N3142);
nor NOR2_1120 (N3325, N3215, N3268);
nor NOR2_1121 (N3326, N3268, N3147);
nor NOR2_1122 (N3327, N3218, N3272);
nor NOR2_1123 (N3328, N3272, N3152);
nor NOR2_1124 (N3329, N3221, N3276);
nor NOR2_1125 (N3330, N3276, N3157);
nor NOR2_1126 (N3331, N3224, N3280);
nor NOR2_1127 (N3332, N3280, N3162);
nor NOR2_1128 (N3333, N3227, N3284);
nor NOR2_1129 (N3334, N3284, N3167);
nor NOR2_1130 (N3335, N3230, N3288);
nor NOR2_1131 (N3336, N3288, N3172);
nor NOR2_1132 (N3337, N3233, N3292);
nor NOR2_1133 (N3338, N3292, N3177);
nor NOR2_1134 (N3339, N3236, N3296);
nor NOR2_1135 (N3340, N3296, N3182);
nor NOR2_1136 (N3341, N3300, N3301);
nor NOR2_1137 (N3344, N3302, N1044);
nor NOR2_1138 (N3348, N3245, N3305);
nor NOR2_1139 (N3349, N3305, N1092);
nor NOR2_1140 (N3350, N3127, N3305);
nor NOR2_1141 (N3353, N3309, N3310);
nor NOR2_1142 (N3356, N3314, N3311);
  nor NOR2_1143 (keyinput_Wire_0[161], N3257, N3317);
  xnor keyGate_0_161(N3360, keyinput161, keyinput_Wire_0[161]);
  nor NOR2_1144 (keyinput_Wire_0[162], N3317, N3254);
  xnor keyGate_0_162(KeyNOTWire_0[82], keyinput162, keyinput_Wire_0[162]);
  not KeyNOTGate_0_82(N3361, KeyNOTWire_0[82]);
  nor NOR2_1145 (keyinput_Wire_0[163], N3321, N3322);
  xnor keyGate_0_163(N3362, keyinput163, keyinput_Wire_0[163]);
nor NOR2_1146 (N3365, N3323, N3324);
nor NOR2_1147 (N3368, N3325, N3326);
nor NOR2_1148 (N3371, N3327, N3328);
nor NOR2_1149 (N3374, N3329, N3330);
nor NOR2_1150 (N3377, N3331, N3332);
nor NOR2_1151 (N3380, N3333, N3334);
nor NOR2_1152 (N3383, N3335, N3336);
nor NOR2_1153 (N3386, N3337, N3338);
nor NOR2_1154 (N3389, N3339, N3340);
nor NOR2_1155 (N3392, N3341, N996);
nor NOR2_1156 (N3396, N3302, N3344);
nor NOR2_1157 (N3397, N3344, N1044);
nor NOR2_1158 (N3398, N3193, N3344);
nor NOR2_1159 (N3401, N3348, N3349);
nor NOR2_1160 (N3404, N3353, N3350);
nor NOR2_1161 (N3408, N3314, N3356);
nor NOR2_1162 (N3409, N3356, N3311);
  nor NOR2_1163 (keyinput_Wire_0[164], N3360, N3361);
  xor keyGate_0_164(KeyNOTWire_0[83], keyinput164, keyinput_Wire_0[164]);
  not KeyNOTGate_0_83(N3410, KeyNOTWire_0[83]);
  nor NOR2_1164 (keyinput_Wire_0[165], N3362, N1239);
  xor keyGate_0_165(KeyNOTWire_0[84], keyinput165, keyinput_Wire_0[165]);
  not KeyNOTGate_0_84(N3413, KeyNOTWire_0[84]);
nor NOR2_1165 (N3417, N3365, N564);
nor NOR2_1166 (N3421, N3368, N612);
nor NOR2_1167 (N3425, N3371, N660);
nor NOR2_1168 (N3429, N3374, N708);
nor NOR2_1169 (N3433, N3377, N756);
nor NOR2_1170 (N3437, N3380, N804);
nor NOR2_1171 (N3441, N3383, N852);
nor NOR2_1172 (N3445, N3386, N900);
nor NOR2_1173 (N3449, N3389, N948);
nor NOR2_1174 (N3453, N3341, N3392);
nor NOR2_1175 (N3454, N3392, N996);
nor NOR2_1176 (N3455, N3239, N3392);
nor NOR2_1177 (N3458, N3396, N3397);
nor NOR2_1178 (N3461, N3401, N3398);
nor NOR2_1179 (N3465, N3353, N3404);
nor NOR2_1180 (N3466, N3404, N3350);
nor NOR2_1181 (N3467, N3408, N3409);
  nor NOR2_1182 (keyinput_Wire_0[166], N3410, N1191);
  xor keyGate_0_166(N3470, keyinput166, keyinput_Wire_0[166]);
  nor NOR2_1183 (keyinput_Wire_0[167], N3362, N3413);
  xor keyGate_0_167(N3474, keyinput167, keyinput_Wire_0[167]);
  nor NOR2_1184 (keyinput_Wire_0[168], N3413, N1239);
  xor keyGate_0_168(KeyNOTWire_0[85], keyinput168, keyinput_Wire_0[168]);
  not KeyNOTGate_0_85(N3475, KeyNOTWire_0[85]);
  nor NOR2_1185 (keyinput_Wire_0[169], N3260, N3413);
  xor keyGate_0_169(KeyNOTWire_0[86], keyinput169, keyinput_Wire_0[169]);
  not KeyNOTGate_0_86(N3476, KeyNOTWire_0[86]);
nor NOR2_1186 (N3479, N3365, N3417);
nor NOR2_1187 (N3480, N3417, N564);
nor NOR2_1188 (N3481, N3264, N3417);
nor NOR2_1189 (N3484, N3368, N3421);
nor NOR2_1190 (N3485, N3421, N612);
nor NOR2_1191 (N3486, N3268, N3421);
nor NOR2_1192 (N3489, N3371, N3425);
nor NOR2_1193 (N3490, N3425, N660);
nor NOR2_1194 (N3491, N3272, N3425);
nor NOR2_1195 (N3494, N3374, N3429);
nor NOR2_1196 (N3495, N3429, N708);
nor NOR2_1197 (N3496, N3276, N3429);
nor NOR2_1198 (N3499, N3377, N3433);
nor NOR2_1199 (N3500, N3433, N756);
nor NOR2_1200 (N3501, N3280, N3433);
nor NOR2_1201 (N3504, N3380, N3437);
nor NOR2_1202 (N3505, N3437, N804);
nor NOR2_1203 (N3506, N3284, N3437);
nor NOR2_1204 (N3509, N3383, N3441);
nor NOR2_1205 (N3510, N3441, N852);
nor NOR2_1206 (N3511, N3288, N3441);
nor NOR2_1207 (N3514, N3386, N3445);
nor NOR2_1208 (N3515, N3445, N900);
nor NOR2_1209 (N3516, N3292, N3445);
nor NOR2_1210 (N3519, N3389, N3449);
nor NOR2_1211 (N3520, N3449, N948);
nor NOR2_1212 (N3521, N3296, N3449);
nor NOR2_1213 (N3524, N3453, N3454);
nor NOR2_1214 (N3527, N3458, N3455);
nor NOR2_1215 (N3531, N3401, N3461);
nor NOR2_1216 (N3532, N3461, N3398);
nor NOR2_1217 (N3533, N3465, N3466);
nor NOR2_1218 (N3536, N3467, N1143);
nor NOR2_1219 (N3540, N3410, N3470);
nor NOR2_1220 (N3541, N3470, N1191);
  nor NOR2_1221 (keyinput_Wire_0[170], N3317, N3470);
  xnor keyGate_0_170(N3542, keyinput170, keyinput_Wire_0[170]);
  nor NOR2_1222 (keyinput_Wire_0[171], N3474, N3475);
  xor keyGate_0_171(N3545, keyinput171, keyinput_Wire_0[171]);
  nor NOR2_1223 (keyinput_Wire_0[172], N1287, N3476);
  xnor keyGate_0_172(KeyNOTWire_0[87], keyinput172, keyinput_Wire_0[172]);
  not KeyNOTGate_0_87(N3548, KeyNOTWire_0[87]);
nor NOR2_1224 (N3552, N3479, N3480);
nor NOR2_1225 (N3553, N3484, N3485);
nor NOR2_1226 (N3556, N3489, N3490);
nor NOR2_1227 (N3559, N3494, N3495);
nor NOR2_1228 (N3562, N3499, N3500);
nor NOR2_1229 (N3565, N3504, N3505);
nor NOR2_1230 (N3568, N3509, N3510);
nor NOR2_1231 (N3571, N3514, N3515);
nor NOR2_1232 (N3574, N3519, N3520);
nor NOR2_1233 (N3577, N3524, N3521);
nor NOR2_1234 (N3581, N3458, N3527);
nor NOR2_1235 (N3582, N3527, N3455);
nor NOR2_1236 (N3583, N3531, N3532);
nor NOR2_1237 (N3586, N3533, N1095);
nor NOR2_1238 (N3590, N3467, N3536);
nor NOR2_1239 (N3591, N3536, N1143);
nor NOR2_1240 (N3592, N3356, N3536);
nor NOR2_1241 (N3595, N3540, N3541);
  nor NOR2_1242 (keyinput_Wire_0[173], N3545, N3542);
  xor keyGate_0_173(KeyNOTWire_0[88], keyinput173, keyinput_Wire_0[173]);
  not KeyNOTGate_0_88(N3598, KeyNOTWire_0[88]);
  nor NOR2_1243 (keyinput_Wire_0[174], N1287, N3548);
  xor keyGate_0_174(KeyNOTWire_0[89], keyinput174, keyinput_Wire_0[174]);
  not KeyNOTGate_0_89(N3602, KeyNOTWire_0[89]);
  nor NOR2_1244 (keyinput_Wire_0[175], N3548, N3476);
  xnor keyGate_0_175(KeyNOTWire_0[90], keyinput175, keyinput_Wire_0[175]);
  not KeyNOTGate_0_90(N3603, KeyNOTWire_0[90]);
nor NOR2_1245 (N3604, N3553, N3481);
nor NOR2_1246 (N3608, N3556, N3486);
nor NOR2_1247 (N3612, N3559, N3491);
nor NOR2_1248 (N3616, N3562, N3496);
nor NOR2_1249 (N3620, N3565, N3501);
nor NOR2_1250 (N3624, N3568, N3506);
nor NOR2_1251 (N3628, N3571, N3511);
nor NOR2_1252 (N3632, N3574, N3516);
nor NOR2_1253 (N3636, N3524, N3577);
  nor NOR2_1254 (keyinput_Wire_0[176], N3577, N3521);
  xnor keyGate_0_176(N3637, keyinput176, keyinput_Wire_0[176]);
nor NOR2_1255 (N3638, N3581, N3582);
nor NOR2_1256 (N3641, N3583, N1047);
nor NOR2_1257 (N3645, N3533, N3586);
nor NOR2_1258 (N3646, N3586, N1095);
nor NOR2_1259 (N3647, N3404, N3586);
nor NOR2_1260 (N3650, N3590, N3591);
nor NOR2_1261 (N3653, N3595, N3592);
  nor NOR2_1262 (keyinput_Wire_0[177], N3545, N3598);
  xnor keyGate_0_177(KeyNOTWire_0[91], keyinput177, keyinput_Wire_0[177]);
  not KeyNOTGate_0_91(N3657, KeyNOTWire_0[91]);
  nor NOR2_1263 (keyinput_Wire_0[178], N3598, N3542);
  xnor keyGate_0_178(N3658, keyinput178, keyinput_Wire_0[178]);
  nor NOR2_1264 (keyinput_Wire_0[179], N3602, N3603);
  xor keyGate_0_179(KeyNOTWire_0[92], keyinput179, keyinput_Wire_0[179]);
  not KeyNOTGate_0_92(N3659, KeyNOTWire_0[92]);
nor NOR2_1265 (N3662, N3553, N3604);
nor NOR2_1266 (N3663, N3604, N3481);
nor NOR2_1267 (N3664, N3556, N3608);
nor NOR2_1268 (N3665, N3608, N3486);
nor NOR2_1269 (N3666, N3559, N3612);
nor NOR2_1270 (N3667, N3612, N3491);
nor NOR2_1271 (N3668, N3562, N3616);
nor NOR2_1272 (N3669, N3616, N3496);
nor NOR2_1273 (N3670, N3565, N3620);
nor NOR2_1274 (N3671, N3620, N3501);
nor NOR2_1275 (N3672, N3568, N3624);
nor NOR2_1276 (N3673, N3624, N3506);
nor NOR2_1277 (N3674, N3571, N3628);
nor NOR2_1278 (N3675, N3628, N3511);
nor NOR2_1279 (N3676, N3574, N3632);
nor NOR2_1280 (N3677, N3632, N3516);
nor NOR2_1281 (N3678, N3636, N3637);
nor NOR2_1282 (N3681, N3638, N999);
nor NOR2_1283 (N3685, N3583, N3641);
nor NOR2_1284 (N3686, N3641, N1047);
nor NOR2_1285 (N3687, N3461, N3641);
nor NOR2_1286 (N3690, N3645, N3646);
nor NOR2_1287 (N3693, N3650, N3647);
nor NOR2_1288 (N3697, N3595, N3653);
nor NOR2_1289 (N3698, N3653, N3592);
  nor NOR2_1290 (keyinput_Wire_0[180], N3657, N3658);
  xor keyGate_0_180(KeyNOTWire_0[93], keyinput180, keyinput_Wire_0[180]);
  not KeyNOTGate_0_93(N3699, KeyNOTWire_0[93]);
  nor NOR2_1291 (keyinput_Wire_0[181], N3659, N1242);
  xor keyGate_0_181(KeyNOTWire_0[94], keyinput181, keyinput_Wire_0[181]);
  not KeyNOTGate_0_94(N3702, KeyNOTWire_0[94]);
nor NOR2_1292 (N3706, N3662, N3663);
nor NOR2_1293 (N3709, N3664, N3665);
nor NOR2_1294 (N3712, N3666, N3667);
nor NOR2_1295 (N3715, N3668, N3669);
nor NOR2_1296 (N3718, N3670, N3671);
nor NOR2_1297 (N3721, N3672, N3673);
nor NOR2_1298 (N3724, N3674, N3675);
nor NOR2_1299 (N3727, N3676, N3677);
nor NOR2_1300 (N3730, N3678, N951);
nor NOR2_1301 (N3734, N3638, N3681);
nor NOR2_1302 (N3735, N3681, N999);
  nor NOR2_1303 (keyinput_Wire_0[182], N3527, N3681);
  xor keyGate_0_182(KeyNOTWire_0[95], keyinput182, keyinput_Wire_0[182]);
  not KeyNOTGate_0_95(N3736, KeyNOTWire_0[95]);
nor NOR2_1304 (N3739, N3685, N3686);
nor NOR2_1305 (N3742, N3690, N3687);
nor NOR2_1306 (N3746, N3650, N3693);
nor NOR2_1307 (N3747, N3693, N3647);
nor NOR2_1308 (N3748, N3697, N3698);
  nor NOR2_1309 (keyinput_Wire_0[183], N3699, N1194);
  xnor keyGate_0_183(KeyNOTWire_0[96], keyinput183, keyinput_Wire_0[183]);
  not KeyNOTGate_0_96(N3751, KeyNOTWire_0[96]);
  nor NOR2_1310 (keyinput_Wire_0[184], N3659, N3702);
  xor keyGate_0_184(KeyNOTWire_0[97], keyinput184, keyinput_Wire_0[184]);
  not KeyNOTGate_0_97(N3755, KeyNOTWire_0[97]);
  nor NOR2_1311 (keyinput_Wire_0[185], N3702, N1242);
  xor keyGate_0_185(KeyNOTWire_0[98], keyinput185, keyinput_Wire_0[185]);
  not KeyNOTGate_0_98(N3756, KeyNOTWire_0[98]);
  nor NOR2_1312 (keyinput_Wire_0[186], N3548, N3702);
  xnor keyGate_0_186(N3757, keyinput186, keyinput_Wire_0[186]);
nor NOR2_1313 (N3760, N3706, N567);
nor NOR2_1314 (N3764, N3709, N615);
nor NOR2_1315 (N3768, N3712, N663);
nor NOR2_1316 (N3772, N3715, N711);
nor NOR2_1317 (N3776, N3718, N759);
nor NOR2_1318 (N3780, N3721, N807);
nor NOR2_1319 (N3784, N3724, N855);
nor NOR2_1320 (N3788, N3727, N903);
nor NOR2_1321 (N3792, N3678, N3730);
nor NOR2_1322 (N3793, N3730, N951);
nor NOR2_1323 (N3794, N3577, N3730);
nor NOR2_1324 (N3797, N3734, N3735);
nor NOR2_1325 (N3800, N3739, N3736);
nor NOR2_1326 (N3804, N3690, N3742);
nor NOR2_1327 (N3805, N3742, N3687);
nor NOR2_1328 (N3806, N3746, N3747);
nor NOR2_1329 (N3809, N3748, N1146);
nor NOR2_1330 (N3813, N3699, N3751);
nor NOR2_1331 (N3814, N3751, N1194);
  nor NOR2_1332 (keyinput_Wire_0[187], N3598, N3751);
  xor keyGate_0_187(N3815, keyinput187, keyinput_Wire_0[187]);
  nor NOR2_1333 (keyinput_Wire_0[188], N3755, N3756);
  xnor keyGate_0_188(N3818, keyinput188, keyinput_Wire_0[188]);
  nor NOR2_1334 (keyinput_Wire_0[189], N1290, N3757);
  xnor keyGate_0_189(KeyNOTWire_0[99], keyinput189, keyinput_Wire_0[189]);
  not KeyNOTGate_0_99(N3821, KeyNOTWire_0[99]);
nor NOR2_1335 (N3825, N3706, N3760);
nor NOR2_1336 (N3826, N3760, N567);
nor NOR2_1337 (N3827, N3604, N3760);
nor NOR2_1338 (N3830, N3709, N3764);
nor NOR2_1339 (N3831, N3764, N615);
nor NOR2_1340 (N3832, N3608, N3764);
nor NOR2_1341 (N3835, N3712, N3768);
nor NOR2_1342 (N3836, N3768, N663);
nor NOR2_1343 (N3837, N3612, N3768);
nor NOR2_1344 (N3840, N3715, N3772);
nor NOR2_1345 (N3841, N3772, N711);
  nor NOR2_1346 (keyinput_Wire_0[190], N3616, N3772);
  xnor keyGate_0_190(KeyNOTWire_0[100], keyinput190, keyinput_Wire_0[190]);
  not KeyNOTGate_0_100(N3842, KeyNOTWire_0[100]);
nor NOR2_1347 (N3845, N3718, N3776);
nor NOR2_1348 (N3846, N3776, N759);
nor NOR2_1349 (N3847, N3620, N3776);
nor NOR2_1350 (N3850, N3721, N3780);
nor NOR2_1351 (N3851, N3780, N807);
nor NOR2_1352 (N3852, N3624, N3780);
nor NOR2_1353 (N3855, N3724, N3784);
nor NOR2_1354 (N3856, N3784, N855);
nor NOR2_1355 (N3857, N3628, N3784);
nor NOR2_1356 (N3860, N3727, N3788);
nor NOR2_1357 (N3861, N3788, N903);
nor NOR2_1358 (N3862, N3632, N3788);
nor NOR2_1359 (N3865, N3792, N3793);
nor NOR2_1360 (N3868, N3797, N3794);
nor NOR2_1361 (N3872, N3739, N3800);
nor NOR2_1362 (N3873, N3800, N3736);
nor NOR2_1363 (N3874, N3804, N3805);
nor NOR2_1364 (N3877, N3806, N1098);
nor NOR2_1365 (N3881, N3748, N3809);
nor NOR2_1366 (N3882, N3809, N1146);
nor NOR2_1367 (N3883, N3653, N3809);
nor NOR2_1368 (N3886, N3813, N3814);
  nor NOR2_1369 (keyinput_Wire_0[191], N3818, N3815);
  xor keyGate_0_191(N3889, keyinput191, keyinput_Wire_0[191]);
  nor NOR2_1370 (keyinput_Wire_0[192], N1290, N3821);
  xnor keyGate_0_192(KeyNOTWire_0[101], keyinput192, keyinput_Wire_0[192]);
  not KeyNOTGate_0_101(N3893, KeyNOTWire_0[101]);
  nor NOR2_1371 (keyinput_Wire_0[193], N3821, N3757);
  xnor keyGate_0_193(KeyNOTWire_0[102], keyinput193, keyinput_Wire_0[193]);
  not KeyNOTGate_0_102(N3894, KeyNOTWire_0[102]);
nor NOR2_1372 (N3895, N3825, N3826);
nor NOR2_1373 (N3896, N3830, N3831);
nor NOR2_1374 (N3899, N3835, N3836);
nor NOR2_1375 (N3902, N3840, N3841);
nor NOR2_1376 (N3905, N3845, N3846);
nor NOR2_1377 (N3908, N3850, N3851);
nor NOR2_1378 (N3911, N3855, N3856);
nor NOR2_1379 (N3914, N3860, N3861);
nor NOR2_1380 (N3917, N3865, N3862);
nor NOR2_1381 (N3921, N3797, N3868);
nor NOR2_1382 (N3922, N3868, N3794);
nor NOR2_1383 (N3923, N3872, N3873);
nor NOR2_1384 (N3926, N3874, N1050);
nor NOR2_1385 (N3930, N3806, N3877);
nor NOR2_1386 (N3931, N3877, N1098);
nor NOR2_1387 (N3932, N3693, N3877);
nor NOR2_1388 (N3935, N3881, N3882);
nor NOR2_1389 (N3938, N3886, N3883);
  nor NOR2_1390 (keyinput_Wire_0[194], N3818, N3889);
  xor keyGate_0_194(KeyNOTWire_0[103], keyinput194, keyinput_Wire_0[194]);
  not KeyNOTGate_0_103(N3942, KeyNOTWire_0[103]);
  nor NOR2_1391 (keyinput_Wire_0[195], N3889, N3815);
  xor keyGate_0_195(KeyNOTWire_0[104], keyinput195, keyinput_Wire_0[195]);
  not KeyNOTGate_0_104(N3943, KeyNOTWire_0[104]);
  nor NOR2_1392 (keyinput_Wire_0[196], N3893, N3894);
  xor keyGate_0_196(KeyNOTWire_0[105], keyinput196, keyinput_Wire_0[196]);
  not KeyNOTGate_0_105(N3944, KeyNOTWire_0[105]);
nor NOR2_1393 (N3947, N3896, N3827);
nor NOR2_1394 (N3951, N3899, N3832);
nor NOR2_1395 (N3955, N3902, N3837);
nor NOR2_1396 (N3959, N3905, N3842);
nor NOR2_1397 (N3963, N3908, N3847);
nor NOR2_1398 (N3967, N3911, N3852);
nor NOR2_1399 (N3971, N3914, N3857);
nor NOR2_1400 (N3975, N3865, N3917);
nor NOR2_1401 (N3976, N3917, N3862);
nor NOR2_1402 (N3977, N3921, N3922);
nor NOR2_1403 (N3980, N3923, N1002);
nor NOR2_1404 (N3984, N3874, N3926);
nor NOR2_1405 (N3985, N3926, N1050);
nor NOR2_1406 (N3986, N3742, N3926);
nor NOR2_1407 (N3989, N3930, N3931);
nor NOR2_1408 (N3992, N3935, N3932);
nor NOR2_1409 (N3996, N3886, N3938);
nor NOR2_1410 (N3997, N3938, N3883);
  nor NOR2_1411 (keyinput_Wire_0[197], N3942, N3943);
  xor keyGate_0_197(KeyNOTWire_0[106], keyinput197, keyinput_Wire_0[197]);
  not KeyNOTGate_0_106(N3998, KeyNOTWire_0[106]);
  nor NOR2_1412 (keyinput_Wire_0[198], N3944, N1245);
  xor keyGate_0_198(N4001, keyinput198, keyinput_Wire_0[198]);
nor NOR2_1413 (N4005, N3896, N3947);
nor NOR2_1414 (N4006, N3947, N3827);
nor NOR2_1415 (N4007, N3899, N3951);
nor NOR2_1416 (N4008, N3951, N3832);
nor NOR2_1417 (N4009, N3902, N3955);
nor NOR2_1418 (N4010, N3955, N3837);
nor NOR2_1419 (N4011, N3905, N3959);
nor NOR2_1420 (N4012, N3959, N3842);
nor NOR2_1421 (N4013, N3908, N3963);
nor NOR2_1422 (N4014, N3963, N3847);
nor NOR2_1423 (N4015, N3911, N3967);
nor NOR2_1424 (N4016, N3967, N3852);
nor NOR2_1425 (N4017, N3914, N3971);
nor NOR2_1426 (N4018, N3971, N3857);
nor NOR2_1427 (N4019, N3975, N3976);
nor NOR2_1428 (N4022, N3977, N954);
nor NOR2_1429 (N4026, N3923, N3980);
nor NOR2_1430 (N4027, N3980, N1002);
nor NOR2_1431 (N4028, N3800, N3980);
nor NOR2_1432 (N4031, N3984, N3985);
nor NOR2_1433 (N4034, N3989, N3986);
nor NOR2_1434 (N4038, N3935, N3992);
nor NOR2_1435 (N4039, N3992, N3932);
nor NOR2_1436 (N4040, N3996, N3997);
  nor NOR2_1437 (keyinput_Wire_0[199], N3998, N1197);
  xor keyGate_0_199(KeyNOTWire_0[107], keyinput199, keyinput_Wire_0[199]);
  not KeyNOTGate_0_107(N4043, KeyNOTWire_0[107]);
  nor NOR2_1438 (keyinput_Wire_0[200], N3944, N4001);
  xor keyGate_0_200(N4047, keyinput200, keyinput_Wire_0[200]);
  nor NOR2_1439 (keyinput_Wire_0[201], N4001, N1245);
  xnor keyGate_0_201(N4048, keyinput201, keyinput_Wire_0[201]);
  nor NOR2_1440 (keyinput_Wire_0[202], N3821, N4001);
  xnor keyGate_0_202(KeyNOTWire_0[108], keyinput202, keyinput_Wire_0[202]);
  not KeyNOTGate_0_108(N4049, KeyNOTWire_0[108]);
nor NOR2_1441 (N4052, N4005, N4006);
nor NOR2_1442 (N4055, N4007, N4008);
nor NOR2_1443 (N4058, N4009, N4010);
nor NOR2_1444 (N4061, N4011, N4012);
nor NOR2_1445 (N4064, N4013, N4014);
nor NOR2_1446 (N4067, N4015, N4016);
nor NOR2_1447 (N4070, N4017, N4018);
nor NOR2_1448 (N4073, N4019, N906);
nor NOR2_1449 (N4077, N3977, N4022);
nor NOR2_1450 (N4078, N4022, N954);
nor NOR2_1451 (N4079, N3868, N4022);
nor NOR2_1452 (N4082, N4026, N4027);
nor NOR2_1453 (N4085, N4031, N4028);
nor NOR2_1454 (N4089, N3989, N4034);
nor NOR2_1455 (N4090, N4034, N3986);
nor NOR2_1456 (N4091, N4038, N4039);
nor NOR2_1457 (N4094, N4040, N1149);
nor NOR2_1458 (N4098, N3998, N4043);
nor NOR2_1459 (N4099, N4043, N1197);
  nor NOR2_1460 (keyinput_Wire_0[203], N3889, N4043);
  xor keyGate_0_203(KeyNOTWire_0[109], keyinput203, keyinput_Wire_0[203]);
  not KeyNOTGate_0_109(N4100, KeyNOTWire_0[109]);
  nor NOR2_1461 (keyinput_Wire_0[204], N4047, N4048);
  xor keyGate_0_204(N4103, keyinput204, keyinput_Wire_0[204]);
  nor NOR2_1462 (keyinput_Wire_0[205], N1293, N4049);
  xor keyGate_0_205(KeyNOTWire_0[110], keyinput205, keyinput_Wire_0[205]);
  not KeyNOTGate_0_110(N4106, KeyNOTWire_0[110]);
nor NOR2_1463 (N4110, N4052, N570);
nor NOR2_1464 (N4114, N4055, N618);
nor NOR2_1465 (N4118, N4058, N666);
nor NOR2_1466 (N4122, N4061, N714);
nor NOR2_1467 (N4126, N4064, N762);
nor NOR2_1468 (N4130, N4067, N810);
nor NOR2_1469 (N4134, N4070, N858);
nor NOR2_1470 (N4138, N4019, N4073);
nor NOR2_1471 (N4139, N4073, N906);
nor NOR2_1472 (N4140, N3917, N4073);
nor NOR2_1473 (N4143, N4077, N4078);
nor NOR2_1474 (N4146, N4082, N4079);
nor NOR2_1475 (N4150, N4031, N4085);
nor NOR2_1476 (N4151, N4085, N4028);
nor NOR2_1477 (N4152, N4089, N4090);
nor NOR2_1478 (N4155, N4091, N1101);
nor NOR2_1479 (N4159, N4040, N4094);
nor NOR2_1480 (N4160, N4094, N1149);
nor NOR2_1481 (N4161, N3938, N4094);
nor NOR2_1482 (N4164, N4098, N4099);
  nor NOR2_1483 (keyinput_Wire_0[206], N4103, N4100);
  xnor keyGate_0_206(KeyNOTWire_0[111], keyinput206, keyinput_Wire_0[206]);
  not KeyNOTGate_0_111(N4167, KeyNOTWire_0[111]);
  nor NOR2_1484 (keyinput_Wire_0[207], N1293, N4106);
  xnor keyGate_0_207(KeyNOTWire_0[112], keyinput207, keyinput_Wire_0[207]);
  not KeyNOTGate_0_112(N4171, KeyNOTWire_0[112]);
  nor NOR2_1485 (keyinput_Wire_0[208], N4106, N4049);
  xnor keyGate_0_208(N4172, keyinput208, keyinput_Wire_0[208]);
nor NOR2_1486 (N4173, N4052, N4110);
nor NOR2_1487 (N4174, N4110, N570);
nor NOR2_1488 (N4175, N3947, N4110);
nor NOR2_1489 (N4178, N4055, N4114);
nor NOR2_1490 (N4179, N4114, N618);
nor NOR2_1491 (N4180, N3951, N4114);
nor NOR2_1492 (N4183, N4058, N4118);
nor NOR2_1493 (N4184, N4118, N666);
nor NOR2_1494 (N4185, N3955, N4118);
nor NOR2_1495 (N4188, N4061, N4122);
nor NOR2_1496 (N4189, N4122, N714);
nor NOR2_1497 (N4190, N3959, N4122);
nor NOR2_1498 (N4193, N4064, N4126);
nor NOR2_1499 (N4194, N4126, N762);
nor NOR2_1500 (N4195, N3963, N4126);
nor NOR2_1501 (N4198, N4067, N4130);
nor NOR2_1502 (N4199, N4130, N810);
nor NOR2_1503 (N4200, N3967, N4130);
nor NOR2_1504 (N4203, N4070, N4134);
nor NOR2_1505 (N4204, N4134, N858);
nor NOR2_1506 (N4205, N3971, N4134);
nor NOR2_1507 (N4208, N4138, N4139);
nor NOR2_1508 (N4211, N4143, N4140);
nor NOR2_1509 (N4215, N4082, N4146);
nor NOR2_1510 (N4216, N4146, N4079);
nor NOR2_1511 (N4217, N4150, N4151);
nor NOR2_1512 (N4220, N4152, N1053);
nor NOR2_1513 (N4224, N4091, N4155);
nor NOR2_1514 (N4225, N4155, N1101);
nor NOR2_1515 (N4226, N3992, N4155);
nor NOR2_1516 (N4229, N4159, N4160);
nor NOR2_1517 (N4232, N4164, N4161);
  nor NOR2_1518 (keyinput_Wire_0[209], N4103, N4167);
  xor keyGate_0_209(N4236, keyinput209, keyinput_Wire_0[209]);
  nor NOR2_1519 (keyinput_Wire_0[210], N4167, N4100);
  xnor keyGate_0_210(KeyNOTWire_0[113], keyinput210, keyinput_Wire_0[210]);
  not KeyNOTGate_0_113(N4237, KeyNOTWire_0[113]);
  nor NOR2_1520 (keyinput_Wire_0[211], N4171, N4172);
  xor keyGate_0_211(KeyNOTWire_0[114], keyinput211, keyinput_Wire_0[211]);
  not KeyNOTGate_0_114(N4238, KeyNOTWire_0[114]);
nor NOR2_1521 (N4241, N4173, N4174);
nor NOR2_1522 (N4242, N4178, N4179);
nor NOR2_1523 (N4245, N4183, N4184);
nor NOR2_1524 (N4248, N4188, N4189);
nor NOR2_1525 (N4251, N4193, N4194);
nor NOR2_1526 (N4254, N4198, N4199);
nor NOR2_1527 (N4257, N4203, N4204);
nor NOR2_1528 (N4260, N4208, N4205);
nor NOR2_1529 (N4264, N4143, N4211);
  nor NOR2_1530 (keyinput_Wire_0[212], N4211, N4140);
  xor keyGate_0_212(N4265, keyinput212, keyinput_Wire_0[212]);
nor NOR2_1531 (N4266, N4215, N4216);
nor NOR2_1532 (N4269, N4217, N1005);
nor NOR2_1533 (N4273, N4152, N4220);
nor NOR2_1534 (N4274, N4220, N1053);
nor NOR2_1535 (N4275, N4034, N4220);
nor NOR2_1536 (N4278, N4224, N4225);
nor NOR2_1537 (N4281, N4229, N4226);
nor NOR2_1538 (N4285, N4164, N4232);
nor NOR2_1539 (N4286, N4232, N4161);
  nor NOR2_1540 (keyinput_Wire_0[213], N4236, N4237);
  xnor keyGate_0_213(KeyNOTWire_0[115], keyinput213, keyinput_Wire_0[213]);
  not KeyNOTGate_0_115(N4287, KeyNOTWire_0[115]);
  nor NOR2_1541 (keyinput_Wire_0[214], N4238, N1248);
  xnor keyGate_0_214(N4290, keyinput214, keyinput_Wire_0[214]);
nor NOR2_1542 (N4294, N4242, N4175);
nor NOR2_1543 (N4298, N4245, N4180);
nor NOR2_1544 (N4302, N4248, N4185);
nor NOR2_1545 (N4306, N4251, N4190);
nor NOR2_1546 (N4310, N4254, N4195);
nor NOR2_1547 (N4314, N4257, N4200);
nor NOR2_1548 (N4318, N4208, N4260);
  nor NOR2_1549 (keyinput_Wire_0[215], N4260, N4205);
  xor keyGate_0_215(KeyNOTWire_0[116], keyinput215, keyinput_Wire_0[215]);
  not KeyNOTGate_0_116(N4319, KeyNOTWire_0[116]);
nor NOR2_1550 (N4320, N4264, N4265);
nor NOR2_1551 (N4323, N4266, N957);
nor NOR2_1552 (N4327, N4217, N4269);
nor NOR2_1553 (N4328, N4269, N1005);
nor NOR2_1554 (N4329, N4085, N4269);
nor NOR2_1555 (N4332, N4273, N4274);
nor NOR2_1556 (N4335, N4278, N4275);
nor NOR2_1557 (N4339, N4229, N4281);
nor NOR2_1558 (N4340, N4281, N4226);
nor NOR2_1559 (N4341, N4285, N4286);
  nor NOR2_1560 (keyinput_Wire_0[216], N4287, N1200);
  xor keyGate_0_216(N4344, keyinput216, keyinput_Wire_0[216]);
  nor NOR2_1561 (keyinput_Wire_0[217], N4238, N4290);
  xnor keyGate_0_217(KeyNOTWire_0[117], keyinput217, keyinput_Wire_0[217]);
  not KeyNOTGate_0_117(N4348, KeyNOTWire_0[117]);
  nor NOR2_1562 (keyinput_Wire_0[218], N4290, N1248);
  xor keyGate_0_218(KeyNOTWire_0[118], keyinput218, keyinput_Wire_0[218]);
  not KeyNOTGate_0_118(N4349, KeyNOTWire_0[118]);
  nor NOR2_1563 (keyinput_Wire_0[219], N4106, N4290);
  xnor keyGate_0_219(N4350, keyinput219, keyinput_Wire_0[219]);
nor NOR2_1564 (N4353, N4242, N4294);
nor NOR2_1565 (N4354, N4294, N4175);
nor NOR2_1566 (N4355, N4245, N4298);
nor NOR2_1567 (N4356, N4298, N4180);
nor NOR2_1568 (N4357, N4248, N4302);
nor NOR2_1569 (N4358, N4302, N4185);
nor NOR2_1570 (N4359, N4251, N4306);
nor NOR2_1571 (N4360, N4306, N4190);
nor NOR2_1572 (N4361, N4254, N4310);
nor NOR2_1573 (N4362, N4310, N4195);
nor NOR2_1574 (N4363, N4257, N4314);
nor NOR2_1575 (N4364, N4314, N4200);
nor NOR2_1576 (N4365, N4318, N4319);
nor NOR2_1577 (N4368, N4320, N909);
nor NOR2_1578 (N4372, N4266, N4323);
nor NOR2_1579 (N4373, N4323, N957);
nor NOR2_1580 (N4374, N4146, N4323);
nor NOR2_1581 (N4377, N4327, N4328);
nor NOR2_1582 (N4380, N4332, N4329);
nor NOR2_1583 (N4384, N4278, N4335);
nor NOR2_1584 (N4385, N4335, N4275);
nor NOR2_1585 (N4386, N4339, N4340);
nor NOR2_1586 (N4389, N4341, N1152);
nor NOR2_1587 (N4393, N4287, N4344);
nor NOR2_1588 (N4394, N4344, N1200);
  nor NOR2_1589 (keyinput_Wire_0[220], N4167, N4344);
  xnor keyGate_0_220(N4395, keyinput220, keyinput_Wire_0[220]);
  nor NOR2_1590 (keyinput_Wire_0[221], N4348, N4349);
  xor keyGate_0_221(N4398, keyinput221, keyinput_Wire_0[221]);
  nor NOR2_1591 (keyinput_Wire_0[222], N1296, N4350);
  xor keyGate_0_222(N4401, keyinput222, keyinput_Wire_0[222]);
nor NOR2_1592 (N4405, N4353, N4354);
nor NOR2_1593 (N4408, N4355, N4356);
nor NOR2_1594 (N4411, N4357, N4358);
  nor NOR2_1595 (keyinput_Wire_0[223], N4359, N4360);
  xor keyGate_0_223(N4414, keyinput223, keyinput_Wire_0[223]);
nor NOR2_1596 (N4417, N4361, N4362);
nor NOR2_1597 (N4420, N4363, N4364);
nor NOR2_1598 (N4423, N4365, N861);
nor NOR2_1599 (N4427, N4320, N4368);
nor NOR2_1600 (N4428, N4368, N909);
nor NOR2_1601 (N4429, N4211, N4368);
nor NOR2_1602 (N4432, N4372, N4373);
nor NOR2_1603 (N4435, N4377, N4374);
nor NOR2_1604 (N4439, N4332, N4380);
nor NOR2_1605 (N4440, N4380, N4329);
nor NOR2_1606 (N4441, N4384, N4385);
nor NOR2_1607 (N4444, N4386, N1104);
nor NOR2_1608 (N4448, N4341, N4389);
nor NOR2_1609 (N4449, N4389, N1152);
nor NOR2_1610 (N4450, N4232, N4389);
nor NOR2_1611 (N4453, N4393, N4394);
  nor NOR2_1612 (keyinput_Wire_0[224], N4398, N4395);
  xor keyGate_0_224(KeyNOTWire_0[119], keyinput224, keyinput_Wire_0[224]);
  not KeyNOTGate_0_119(N4456, KeyNOTWire_0[119]);
  nor NOR2_1613 (keyinput_Wire_0[225], N1296, N4401);
  xnor keyGate_0_225(KeyNOTWire_0[120], keyinput225, keyinput_Wire_0[225]);
  not KeyNOTGate_0_120(N4460, KeyNOTWire_0[120]);
  nor NOR2_1614 (keyinput_Wire_0[226], N4401, N4350);
  xnor keyGate_0_226(N4461, keyinput226, keyinput_Wire_0[226]);
nor NOR2_1615 (N4462, N4405, N573);
nor NOR2_1616 (N4466, N4408, N621);
  nor NOR2_1617 (keyinput_Wire_0[227], N4411, N669);
  xnor keyGate_0_227(KeyNOTWire_0[121], keyinput227, keyinput_Wire_0[227]);
  not KeyNOTGate_0_121(N4470, KeyNOTWire_0[121]);
nor NOR2_1618 (N4474, N4414, N717);
nor NOR2_1619 (N4478, N4417, N765);
nor NOR2_1620 (N4482, N4420, N813);
nor NOR2_1621 (N4486, N4365, N4423);
nor NOR2_1622 (N4487, N4423, N861);
nor NOR2_1623 (N4488, N4260, N4423);
nor NOR2_1624 (N4491, N4427, N4428);
nor NOR2_1625 (N4494, N4432, N4429);
nor NOR2_1626 (N4498, N4377, N4435);
nor NOR2_1627 (N4499, N4435, N4374);
nor NOR2_1628 (N4500, N4439, N4440);
nor NOR2_1629 (N4503, N4441, N1056);
nor NOR2_1630 (N4507, N4386, N4444);
nor NOR2_1631 (N4508, N4444, N1104);
nor NOR2_1632 (N4509, N4281, N4444);
nor NOR2_1633 (N4512, N4448, N4449);
nor NOR2_1634 (N4515, N4453, N4450);
  nor NOR2_1635 (keyinput_Wire_0[228], N4398, N4456);
  xnor keyGate_0_228(N4519, keyinput228, keyinput_Wire_0[228]);
  nor NOR2_1636 (keyinput_Wire_0[229], N4456, N4395);
  xor keyGate_0_229(KeyNOTWire_0[122], keyinput229, keyinput_Wire_0[229]);
  not KeyNOTGate_0_122(N4520, KeyNOTWire_0[122]);
  nor NOR2_1637 (keyinput_Wire_0[230], N4460, N4461);
  xnor keyGate_0_230(N4521, keyinput230, keyinput_Wire_0[230]);
nor NOR2_1638 (N4524, N4405, N4462);
nor NOR2_1639 (N4525, N4462, N573);
nor NOR2_1640 (N4526, N4294, N4462);
nor NOR2_1641 (N4529, N4408, N4466);
nor NOR2_1642 (N4530, N4466, N621);
nor NOR2_1643 (N4531, N4298, N4466);
nor NOR2_1644 (N4534, N4411, N4470);
nor NOR2_1645 (N4535, N4470, N669);
nor NOR2_1646 (N4536, N4302, N4470);
nor NOR2_1647 (N4539, N4414, N4474);
nor NOR2_1648 (N4540, N4474, N717);
nor NOR2_1649 (N4541, N4306, N4474);
nor NOR2_1650 (N4544, N4417, N4478);
nor NOR2_1651 (N4545, N4478, N765);
nor NOR2_1652 (N4546, N4310, N4478);
nor NOR2_1653 (N4549, N4420, N4482);
nor NOR2_1654 (N4550, N4482, N813);
nor NOR2_1655 (N4551, N4314, N4482);
nor NOR2_1656 (N4554, N4486, N4487);
nor NOR2_1657 (N4557, N4491, N4488);
nor NOR2_1658 (N4561, N4432, N4494);
nor NOR2_1659 (N4562, N4494, N4429);
nor NOR2_1660 (N4563, N4498, N4499);
nor NOR2_1661 (N4566, N4500, N1008);
nor NOR2_1662 (N4570, N4441, N4503);
nor NOR2_1663 (N4571, N4503, N1056);
nor NOR2_1664 (N4572, N4335, N4503);
nor NOR2_1665 (N4575, N4507, N4508);
nor NOR2_1666 (N4578, N4512, N4509);
nor NOR2_1667 (N4582, N4453, N4515);
nor NOR2_1668 (N4583, N4515, N4450);
  nor NOR2_1669 (keyinput_Wire_0[231], N4519, N4520);
  xor keyGate_0_231(KeyNOTWire_0[123], keyinput231, keyinput_Wire_0[231]);
  not KeyNOTGate_0_123(N4584, KeyNOTWire_0[123]);
  nor NOR2_1670 (keyinput_Wire_0[232], N4521, N1251);
  xor keyGate_0_232(N4587, keyinput232, keyinput_Wire_0[232]);
nor NOR2_1671 (N4591, N4524, N4525);
nor NOR2_1672 (N4592, N4529, N4530);
nor NOR2_1673 (N4595, N4534, N4535);
nor NOR2_1674 (N4598, N4539, N4540);
nor NOR2_1675 (N4601, N4544, N4545);
nor NOR2_1676 (N4604, N4549, N4550);
nor NOR2_1677 (N4607, N4554, N4551);
nor NOR2_1678 (N4611, N4491, N4557);
nor NOR2_1679 (N4612, N4557, N4488);
nor NOR2_1680 (N4613, N4561, N4562);
nor NOR2_1681 (N4616, N4563, N960);
nor NOR2_1682 (N4620, N4500, N4566);
nor NOR2_1683 (N4621, N4566, N1008);
nor NOR2_1684 (N4622, N4380, N4566);
nor NOR2_1685 (N4625, N4570, N4571);
nor NOR2_1686 (N4628, N4575, N4572);
nor NOR2_1687 (N4632, N4512, N4578);
nor NOR2_1688 (N4633, N4578, N4509);
nor NOR2_1689 (N4634, N4582, N4583);
  nor NOR2_1690 (keyinput_Wire_0[233], N4584, N1203);
  xor keyGate_0_233(KeyNOTWire_0[124], keyinput233, keyinput_Wire_0[233]);
  not KeyNOTGate_0_124(N4637, KeyNOTWire_0[124]);
  nor NOR2_1691 (keyinput_Wire_0[234], N4521, N4587);
  xor keyGate_0_234(KeyNOTWire_0[125], keyinput234, keyinput_Wire_0[234]);
  not KeyNOTGate_0_125(N4641, KeyNOTWire_0[125]);
  nor NOR2_1692 (keyinput_Wire_0[235], N4587, N1251);
  xor keyGate_0_235(KeyNOTWire_0[126], keyinput235, keyinput_Wire_0[235]);
  not KeyNOTGate_0_126(N4642, KeyNOTWire_0[126]);
nor NOR2_1693 (N4643, N4401, N4587);
nor NOR2_1694 (N4646, N4592, N4526);
nor NOR2_1695 (N4650, N4595, N4531);
nor NOR2_1696 (N4654, N4598, N4536);
nor NOR2_1697 (N4658, N4601, N4541);
nor NOR2_1698 (N4662, N4604, N4546);
nor NOR2_1699 (N4666, N4554, N4607);
nor NOR2_1700 (N4667, N4607, N4551);
nor NOR2_1701 (N4668, N4611, N4612);
nor NOR2_1702 (N4671, N4613, N912);
nor NOR2_1703 (N4675, N4563, N4616);
nor NOR2_1704 (N4676, N4616, N960);
nor NOR2_1705 (N4677, N4435, N4616);
nor NOR2_1706 (N4680, N4620, N4621);
nor NOR2_1707 (N4683, N4625, N4622);
nor NOR2_1708 (N4687, N4575, N4628);
nor NOR2_1709 (N4688, N4628, N4572);
nor NOR2_1710 (N4689, N4632, N4633);
nor NOR2_1711 (N4692, N4634, N1155);
nor NOR2_1712 (N4696, N4584, N4637);
nor NOR2_1713 (N4697, N4637, N1203);
  nor NOR2_1714 (keyinput_Wire_0[236], N4456, N4637);
  xor keyGate_0_236(N4698, keyinput236, keyinput_Wire_0[236]);
  nor NOR2_1715 (keyinput_Wire_0[237], N4641, N4642);
  xnor keyGate_0_237(KeyNOTWire_0[127], keyinput237, keyinput_Wire_0[237]);
  not KeyNOTGate_0_127(N4701, KeyNOTWire_0[127]);
nor NOR2_1716 (N4704, N1299, N4643);
nor NOR2_1717 (N4708, N4592, N4646);
nor NOR2_1718 (N4709, N4646, N4526);
nor NOR2_1719 (N4710, N4595, N4650);
nor NOR2_1720 (N4711, N4650, N4531);
nor NOR2_1721 (N4712, N4598, N4654);
nor NOR2_1722 (N4713, N4654, N4536);
nor NOR2_1723 (N4714, N4601, N4658);
nor NOR2_1724 (N4715, N4658, N4541);
nor NOR2_1725 (N4716, N4604, N4662);
nor NOR2_1726 (N4717, N4662, N4546);
nor NOR2_1727 (N4718, N4666, N4667);
nor NOR2_1728 (N4721, N4668, N864);
nor NOR2_1729 (N4725, N4613, N4671);
nor NOR2_1730 (N4726, N4671, N912);
nor NOR2_1731 (N4727, N4494, N4671);
nor NOR2_1732 (N4730, N4675, N4676);
nor NOR2_1733 (N4733, N4680, N4677);
nor NOR2_1734 (N4737, N4625, N4683);
nor NOR2_1735 (N4738, N4683, N4622);
nor NOR2_1736 (N4739, N4687, N4688);
nor NOR2_1737 (N4742, N4689, N1107);
nor NOR2_1738 (N4746, N4634, N4692);
nor NOR2_1739 (N4747, N4692, N1155);
nor NOR2_1740 (N4748, N4515, N4692);
nor NOR2_1741 (N4751, N4696, N4697);
  nor NOR2_1742 (keyinput_Wire_0[238], N4701, N4698);
  xor keyGate_0_238(KeyNOTWire_0[128], keyinput238, keyinput_Wire_0[238]);
  not KeyNOTGate_0_128(N4754, KeyNOTWire_0[128]);
  nor NOR2_1743 (keyinput_Wire_0[239], N1299, N4704);
  xor keyGate_0_239(N4758, keyinput239, keyinput_Wire_0[239]);
nor NOR2_1744 (N4759, N4704, N4643);
nor NOR2_1745 (N4760, N4708, N4709);
nor NOR2_1746 (N4763, N4710, N4711);
nor NOR2_1747 (N4766, N4712, N4713);
nor NOR2_1748 (N4769, N4714, N4715);
  nor NOR2_1749 (keyinput_Wire_0[240], N4716, N4717);
  xnor keyGate_0_240(KeyNOTWire_0[129], keyinput240, keyinput_Wire_0[240]);
  not KeyNOTGate_0_129(N4772, KeyNOTWire_0[129]);
nor NOR2_1750 (N4775, N4718, N816);
nor NOR2_1751 (N4779, N4668, N4721);
nor NOR2_1752 (N4780, N4721, N864);
nor NOR2_1753 (N4781, N4557, N4721);
nor NOR2_1754 (N4784, N4725, N4726);
nor NOR2_1755 (N4787, N4730, N4727);
nor NOR2_1756 (N4791, N4680, N4733);
nor NOR2_1757 (N4792, N4733, N4677);
nor NOR2_1758 (N4793, N4737, N4738);
nor NOR2_1759 (N4796, N4739, N1059);
nor NOR2_1760 (N4800, N4689, N4742);
nor NOR2_1761 (N4801, N4742, N1107);
nor NOR2_1762 (N4802, N4578, N4742);
nor NOR2_1763 (N4805, N4746, N4747);
nor NOR2_1764 (N4808, N4751, N4748);
  nor NOR2_1765 (keyinput_Wire_0[241], N4701, N4754);
  xor keyGate_0_241(KeyNOTWire_0[130], keyinput241, keyinput_Wire_0[241]);
  not KeyNOTGate_0_130(N4812, KeyNOTWire_0[130]);
  nor NOR2_1766 (keyinput_Wire_0[242], N4754, N4698);
  xnor keyGate_0_242(KeyNOTWire_0[131], keyinput242, keyinput_Wire_0[242]);
  not KeyNOTGate_0_131(N4813, KeyNOTWire_0[131]);
nor NOR2_1767 (N4814, N4758, N4759);
nor NOR2_1768 (N4817, N4760, N576);
nor NOR2_1769 (N4821, N4763, N624);
nor NOR2_1770 (N4825, N4766, N672);
nor NOR2_1771 (N4829, N4769, N720);
nor NOR2_1772 (N4833, N4772, N768);
nor NOR2_1773 (N4837, N4718, N4775);
nor NOR2_1774 (N4838, N4775, N816);
nor NOR2_1775 (N4839, N4607, N4775);
nor NOR2_1776 (N4842, N4779, N4780);
nor NOR2_1777 (N4845, N4784, N4781);
nor NOR2_1778 (N4849, N4730, N4787);
nor NOR2_1779 (N4850, N4787, N4727);
nor NOR2_1780 (N4851, N4791, N4792);
nor NOR2_1781 (N4854, N4793, N1011);
nor NOR2_1782 (N4858, N4739, N4796);
nor NOR2_1783 (N4859, N4796, N1059);
nor NOR2_1784 (N4860, N4628, N4796);
nor NOR2_1785 (N4863, N4800, N4801);
nor NOR2_1786 (N4866, N4805, N4802);
nor NOR2_1787 (N4870, N4751, N4808);
nor NOR2_1788 (N4871, N4808, N4748);
  nor NOR2_1789 (keyinput_Wire_0[243], N4812, N4813);
  xnor keyGate_0_243(KeyNOTWire_0[132], keyinput243, keyinput_Wire_0[243]);
  not KeyNOTGate_0_132(N4872, KeyNOTWire_0[132]);
nor NOR2_1790 (N4875, N4814, N1254);
nor NOR2_1791 (N4879, N4760, N4817);
nor NOR2_1792 (N4880, N4817, N576);
nor NOR2_1793 (N4881, N4646, N4817);
nor NOR2_1794 (N4884, N4763, N4821);
nor NOR2_1795 (N4885, N4821, N624);
nor NOR2_1796 (N4886, N4650, N4821);
nor NOR2_1797 (N4889, N4766, N4825);
nor NOR2_1798 (N4890, N4825, N672);
nor NOR2_1799 (N4891, N4654, N4825);
nor NOR2_1800 (N4894, N4769, N4829);
nor NOR2_1801 (N4895, N4829, N720);
nor NOR2_1802 (N4896, N4658, N4829);
nor NOR2_1803 (N4899, N4772, N4833);
nor NOR2_1804 (N4900, N4833, N768);
nor NOR2_1805 (N4901, N4662, N4833);
nor NOR2_1806 (N4904, N4837, N4838);
nor NOR2_1807 (N4907, N4842, N4839);
nor NOR2_1808 (N4911, N4784, N4845);
nor NOR2_1809 (N4912, N4845, N4781);
nor NOR2_1810 (N4913, N4849, N4850);
nor NOR2_1811 (N4916, N4851, N963);
nor NOR2_1812 (N4920, N4793, N4854);
nor NOR2_1813 (N4921, N4854, N1011);
nor NOR2_1814 (N4922, N4683, N4854);
nor NOR2_1815 (N4925, N4858, N4859);
nor NOR2_1816 (N4928, N4863, N4860);
nor NOR2_1817 (N4932, N4805, N4866);
nor NOR2_1818 (N4933, N4866, N4802);
nor NOR2_1819 (N4934, N4870, N4871);
  nor NOR2_1820 (keyinput_Wire_0[244], N4872, N1206);
  xor keyGate_0_244(KeyNOTWire_0[133], keyinput244, keyinput_Wire_0[244]);
  not KeyNOTGate_0_133(N4937, KeyNOTWire_0[133]);
  nor NOR2_1821 (keyinput_Wire_0[245], N4814, N4875);
  xnor keyGate_0_245(KeyNOTWire_0[134], keyinput245, keyinput_Wire_0[245]);
  not KeyNOTGate_0_134(N4941, KeyNOTWire_0[134]);
nor NOR2_1822 (N4942, N4875, N1254);
nor NOR2_1823 (N4943, N4704, N4875);
nor NOR2_1824 (KeyWire_0_1, N4879, N4880);
  xor flip_it (N4946, KeyWire_0_1, KeyWire_0_2 );
nor NOR2_1825 (N4947, N4884, N4885);
nor NOR2_1826 (N4950, N4889, N4890);
nor NOR2_1827 (N4953, N4894, N4895);
nor NOR2_1828 (N4956, N4899, N4900);
nor NOR2_1829 (N4959, N4904, N4901);
nor NOR2_1830 (N4963, N4842, N4907);
nor NOR2_1831 (N4964, N4907, N4839);
nor NOR2_1832 (N4965, N4911, N4912);
nor NOR2_1833 (N4968, N4913, N915);
nor NOR2_1834 (N4972, N4851, N4916);
nor NOR2_1835 (N4973, N4916, N963);
nor NOR2_1836 (N4974, N4733, N4916);
nor NOR2_1837 (N4977, N4920, N4921);
nor NOR2_1838 (N4980, N4925, N4922);
nor NOR2_1839 (N4984, N4863, N4928);
nor NOR2_1840 (N4985, N4928, N4860);
nor NOR2_1841 (N4986, N4932, N4933);
nor NOR2_1842 (N4989, N4934, N1158);
nor NOR2_1843 (N4993, N4872, N4937);
nor NOR2_1844 (N4994, N4937, N1206);
nor NOR2_1845 (N4995, N4754, N4937);
nor NOR2_1846 (N4998, N4941, N4942);
nor NOR2_1847 (N5001, N1302, N4943);
nor NOR2_1848 (N5005, N4947, N4881);
nor NOR2_1849 (N5009, N4950, N4886);
nor NOR2_1850 (N5013, N4953, N4891);
nor NOR2_1851 (N5017, N4956, N4896);
nor NOR2_1852 (N5021, N4904, N4959);
nor NOR2_1853 (N5022, N4959, N4901);
nor NOR2_1854 (N5023, N4963, N4964);
nor NOR2_1855 (N5026, N4965, N867);
nor NOR2_1856 (N5030, N4913, N4968);
nor NOR2_1857 (N5031, N4968, N915);
nor NOR2_1858 (N5032, N4787, N4968);
nor NOR2_1859 (N5035, N4972, N4973);
nor NOR2_1860 (N5038, N4977, N4974);
nor NOR2_1861 (N5042, N4925, N4980);
nor NOR2_1862 (N5043, N4980, N4922);
nor NOR2_1863 (N5044, N4984, N4985);
nor NOR2_1864 (N5047, N4986, N1110);
nor NOR2_1865 (N5051, N4934, N4989);
nor NOR2_1866 (N5052, N4989, N1158);
nor NOR2_1867 (N5053, N4808, N4989);
nor NOR2_1868 (N5056, N4993, N4994);
  nor NOR2_1869 (keyinput_Wire_0[246], N4998, N4995);
  xor keyGate_0_246(N5059, keyinput246, keyinput_Wire_0[246]);
nor NOR2_1870 (N5063, N1302, N5001);
nor NOR2_1871 (N5064, N5001, N4943);
nor NOR2_1872 (N5065, N4947, N5005);
nor NOR2_1873 (N5066, N5005, N4881);
nor NOR2_1874 (N5067, N4950, N5009);
nor NOR2_1875 (N5068, N5009, N4886);
nor NOR2_1876 (N5069, N4953, N5013);
nor NOR2_1877 (N5070, N5013, N4891);
nor NOR2_1878 (N5071, N4956, N5017);
nor NOR2_1879 (N5072, N5017, N4896);
nor NOR2_1880 (N5073, N5021, N5022);
nor NOR2_1881 (N5076, N5023, N819);
nor NOR2_1882 (N5080, N4965, N5026);
nor NOR2_1883 (N5081, N5026, N867);
nor NOR2_1884 (N5082, N4845, N5026);
nor NOR2_1885 (N5085, N5030, N5031);
nor NOR2_1886 (N5088, N5035, N5032);
nor NOR2_1887 (N5092, N4977, N5038);
nor NOR2_1888 (N5093, N5038, N4974);
nor NOR2_1889 (N5094, N5042, N5043);
nor NOR2_1890 (N5097, N5044, N1062);
nor NOR2_1891 (N5101, N4986, N5047);
nor NOR2_1892 (N5102, N5047, N1110);
nor NOR2_1893 (N5103, N4866, N5047);
nor NOR2_1894 (N5106, N5051, N5052);
nor NOR2_1895 (N5109, N5056, N5053);
nor NOR2_1896 (N5113, N4998, N5059);
  nor NOR2_1897 (keyinput_Wire_0[247], N5059, N4995);
  xnor keyGate_0_247(KeyNOTWire_0[135], keyinput247, keyinput_Wire_0[247]);
  not KeyNOTGate_0_135(N5114, KeyNOTWire_0[135]);
nor NOR2_1898 (N5115, N5063, N5064);
nor NOR2_1899 (N5118, N5065, N5066);
nor NOR2_1900 (N5121, N5067, N5068);
nor NOR2_1901 (N5124, N5069, N5070);
nor NOR2_1902 (N5127, N5071, N5072);
nor NOR2_1903 (N5130, N5073, N771);
nor NOR2_1904 (N5134, N5023, N5076);
nor NOR2_1905 (N5135, N5076, N819);
nor NOR2_1906 (N5136, N4907, N5076);
nor NOR2_1907 (N5139, N5080, N5081);
nor NOR2_1908 (N5142, N5085, N5082);
nor NOR2_1909 (N5146, N5035, N5088);
nor NOR2_1910 (N5147, N5088, N5032);
nor NOR2_1911 (N5148, N5092, N5093);
nor NOR2_1912 (N5151, N5094, N1014);
nor NOR2_1913 (N5155, N5044, N5097);
nor NOR2_1914 (N5156, N5097, N1062);
nor NOR2_1915 (N5157, N4928, N5097);
nor NOR2_1916 (N5160, N5101, N5102);
nor NOR2_1917 (N5163, N5106, N5103);
nor NOR2_1918 (N5167, N5056, N5109);
nor NOR2_1919 (N5168, N5109, N5053);
  nor NOR2_1920 (keyinput_Wire_0[248], N5113, N5114);
  xor keyGate_0_248(N5169, keyinput248, keyinput_Wire_0[248]);
nor NOR2_1921 (N5172, N5115, N1257);
nor NOR2_1922 (N5176, N5118, N579);
nor NOR2_1923 (N5180, N5121, N627);
nor NOR2_1924 (N5184, N5124, N675);
nor NOR2_1925 (N5188, N5127, N723);
nor NOR2_1926 (N5192, N5073, N5130);
nor NOR2_1927 (N5193, N5130, N771);
nor NOR2_1928 (N5194, N4959, N5130);
nor NOR2_1929 (N5197, N5134, N5135);
nor NOR2_1930 (N5200, N5139, N5136);
nor NOR2_1931 (N5204, N5085, N5142);
nor NOR2_1932 (N5205, N5142, N5082);
nor NOR2_1933 (N5206, N5146, N5147);
nor NOR2_1934 (N5209, N5148, N966);
nor NOR2_1935 (N5213, N5094, N5151);
nor NOR2_1936 (N5214, N5151, N1014);
nor NOR2_1937 (N5215, N4980, N5151);
nor NOR2_1938 (N5218, N5155, N5156);
nor NOR2_1939 (N5221, N5160, N5157);
nor NOR2_1940 (N5225, N5106, N5163);
nor NOR2_1941 (N5226, N5163, N5103);
nor NOR2_1942 (N5227, N5167, N5168);
  nor NOR2_1943 (keyinput_Wire_0[249], N5169, N1209);
  xnor keyGate_0_249(KeyNOTWire_0[136], keyinput249, keyinput_Wire_0[249]);
  not KeyNOTGate_0_136(N5230, KeyNOTWire_0[136]);
nor NOR2_1944 (N5234, N5115, N5172);
nor NOR2_1945 (N5235, N5172, N1257);
nor NOR2_1946 (N5236, N5001, N5172);
nor NOR2_1947 (N5239, N5118, N5176);
nor NOR2_1948 (N5240, N5176, N579);
nor NOR2_1949 (N5241, N5005, N5176);
nor NOR2_1950 (N5244, N5121, N5180);
nor NOR2_1951 (N5245, N5180, N627);
nor NOR2_1952 (N5246, N5009, N5180);
nor NOR2_1953 (N5249, N5124, N5184);
nor NOR2_1954 (N5250, N5184, N675);
nor NOR2_1955 (N5251, N5013, N5184);
nor NOR2_1956 (N5254, N5127, N5188);
nor NOR2_1957 (N5255, N5188, N723);
nor NOR2_1958 (N5256, N5017, N5188);
nor NOR2_1959 (N5259, N5192, N5193);
nor NOR2_1960 (N5262, N5197, N5194);
nor NOR2_1961 (N5266, N5139, N5200);
nor NOR2_1962 (N5267, N5200, N5136);
nor NOR2_1963 (N5268, N5204, N5205);
nor NOR2_1964 (N5271, N5206, N918);
nor NOR2_1965 (N5275, N5148, N5209);
nor NOR2_1966 (N5276, N5209, N966);
nor NOR2_1967 (N5277, N5038, N5209);
nor NOR2_1968 (N5280, N5213, N5214);
nor NOR2_1969 (N5283, N5218, N5215);
nor NOR2_1970 (N5287, N5160, N5221);
nor NOR2_1971 (N5288, N5221, N5157);
nor NOR2_1972 (N5289, N5225, N5226);
nor NOR2_1973 (N5292, N5227, N1161);
nor NOR2_1974 (N5296, N5169, N5230);
nor NOR2_1975 (N5297, N5230, N1209);
  nor NOR2_1976 (keyinput_Wire_0[250], N5059, N5230);
  xnor keyGate_0_250(KeyNOTWire_0[137], keyinput250, keyinput_Wire_0[250]);
  not KeyNOTGate_0_137(N5298, KeyNOTWire_0[137]);
nor NOR2_1977 (N5301, N5234, N5235);
nor NOR2_1978 (N5304, N1305, N5236);
nor NOR2_1979 (N5308, N5239, N5240);
nor NOR2_1980 (N5309, N5244, N5245);
nor NOR2_1981 (N5312, N5249, N5250);
nor NOR2_1982 (N5315, N5254, N5255);
nor NOR2_1983 (N5318, N5259, N5256);
nor NOR2_1984 (N5322, N5197, N5262);
nor NOR2_1985 (N5323, N5262, N5194);
nor NOR2_1986 (N5324, N5266, N5267);
nor NOR2_1987 (N5327, N5268, N870);
nor NOR2_1988 (N5331, N5206, N5271);
nor NOR2_1989 (N5332, N5271, N918);
nor NOR2_1990 (N5333, N5088, N5271);
nor NOR2_1991 (N5336, N5275, N5276);
nor NOR2_1992 (N5339, N5280, N5277);
nor NOR2_1993 (N5343, N5218, N5283);
nor NOR2_1994 (N5344, N5283, N5215);
nor NOR2_1995 (N5345, N5287, N5288);
nor NOR2_1996 (N5348, N5289, N1113);
nor NOR2_1997 (N5352, N5227, N5292);
nor NOR2_1998 (N5353, N5292, N1161);
nor NOR2_1999 (N5354, N5109, N5292);
nor NOR2_2000 (N5357, N5296, N5297);
nor NOR2_2001 (N5360, N5301, N5298);
nor NOR2_2002 (N5364, N1305, N5304);
nor NOR2_2003 (N5365, N5304, N5236);
nor NOR2_2004 (N5366, N5309, N5241);
nor NOR2_2005 (N5370, N5312, N5246);
nor NOR2_2006 (N5374, N5315, N5251);
nor NOR2_2007 (N5378, N5259, N5318);
nor NOR2_2008 (N5379, N5318, N5256);
nor NOR2_2009 (N5380, N5322, N5323);
nor NOR2_2010 (N5383, N5324, N822);
nor NOR2_2011 (N5387, N5268, N5327);
nor NOR2_2012 (N5388, N5327, N870);
nor NOR2_2013 (N5389, N5142, N5327);
nor NOR2_2014 (N5392, N5331, N5332);
nor NOR2_2015 (N5395, N5336, N5333);
nor NOR2_2016 (N5399, N5280, N5339);
nor NOR2_2017 (N5400, N5339, N5277);
nor NOR2_2018 (N5401, N5343, N5344);
nor NOR2_2019 (N5404, N5345, N1065);
nor NOR2_2020 (N5408, N5289, N5348);
nor NOR2_2021 (N5409, N5348, N1113);
nor NOR2_2022 (N5410, N5163, N5348);
nor NOR2_2023 (N5413, N5352, N5353);
nor NOR2_2024 (N5416, N5357, N5354);
  nor NOR2_2025 (keyinput_Wire_0[251], N5301, N5360);
  xor keyGate_0_251(KeyNOTWire_0[138], keyinput251, keyinput_Wire_0[251]);
  not KeyNOTGate_0_138(N5420, KeyNOTWire_0[138]);
nor NOR2_2026 (N5421, N5360, N5298);
nor NOR2_2027 (N5422, N5364, N5365);
nor NOR2_2028 (N5425, N5309, N5366);
nor NOR2_2029 (N5426, N5366, N5241);
nor NOR2_2030 (N5427, N5312, N5370);
nor NOR2_2031 (N5428, N5370, N5246);
nor NOR2_2032 (N5429, N5315, N5374);
nor NOR2_2033 (N5430, N5374, N5251);
nor NOR2_2034 (N5431, N5378, N5379);
nor NOR2_2035 (N5434, N5380, N774);
nor NOR2_2036 (N5438, N5324, N5383);
nor NOR2_2037 (N5439, N5383, N822);
nor NOR2_2038 (N5440, N5200, N5383);
nor NOR2_2039 (N5443, N5387, N5388);
nor NOR2_2040 (N5446, N5392, N5389);
nor NOR2_2041 (N5450, N5336, N5395);
nor NOR2_2042 (N5451, N5395, N5333);
nor NOR2_2043 (N5452, N5399, N5400);
nor NOR2_2044 (N5455, N5401, N1017);
nor NOR2_2045 (N5459, N5345, N5404);
nor NOR2_2046 (N5460, N5404, N1065);
nor NOR2_2047 (N5461, N5221, N5404);
nor NOR2_2048 (N5464, N5408, N5409);
nor NOR2_2049 (N5467, N5413, N5410);
nor NOR2_2050 (N5471, N5357, N5416);
nor NOR2_2051 (N5472, N5416, N5354);
nor NOR2_2052 (N5473, N5420, N5421);
nor NOR2_2053 (N5476, N5422, N1260);
nor NOR2_2054 (N5480, N5425, N5426);
nor NOR2_2055 (N5483, N5427, N5428);
nor NOR2_2056 (N5486, N5429, N5430);
nor NOR2_2057 (N5489, N5431, N726);
nor NOR2_2058 (N5493, N5380, N5434);
nor NOR2_2059 (N5494, N5434, N774);
nor NOR2_2060 (N5495, N5262, N5434);
nor NOR2_2061 (N5498, N5438, N5439);
nor NOR2_2062 (N5501, N5443, N5440);
nor NOR2_2063 (N5505, N5392, N5446);
nor NOR2_2064 (N5506, N5446, N5389);
nor NOR2_2065 (N5507, N5450, N5451);
nor NOR2_2066 (N5510, N5452, N969);
nor NOR2_2067 (N5514, N5401, N5455);
nor NOR2_2068 (N5515, N5455, N1017);
nor NOR2_2069 (N5516, N5283, N5455);
nor NOR2_2070 (N5519, N5459, N5460);
nor NOR2_2071 (N5522, N5464, N5461);
nor NOR2_2072 (N5526, N5413, N5467);
nor NOR2_2073 (N5527, N5467, N5410);
nor NOR2_2074 (N5528, N5471, N5472);
nor NOR2_2075 (N5531, N5473, N1212);
nor NOR2_2076 (N5535, N5422, N5476);
nor NOR2_2077 (N5536, N5476, N1260);
nor NOR2_2078 (N5537, N5304, N5476);
nor NOR2_2079 (N5540, N5480, N582);
nor NOR2_2080 (N5544, N5483, N630);
nor NOR2_2081 (N5548, N5486, N678);
nor NOR2_2082 (N5552, N5431, N5489);
nor NOR2_2083 (N5553, N5489, N726);
nor NOR2_2084 (N5554, N5318, N5489);
nor NOR2_2085 (N5557, N5493, N5494);
nor NOR2_2086 (N5560, N5498, N5495);
nor NOR2_2087 (N5564, N5443, N5501);
nor NOR2_2088 (N5565, N5501, N5440);
nor NOR2_2089 (N5566, N5505, N5506);
nor NOR2_2090 (N5569, N5507, N921);
nor NOR2_2091 (N5573, N5452, N5510);
nor NOR2_2092 (N5574, N5510, N969);
nor NOR2_2093 (N5575, N5339, N5510);
nor NOR2_2094 (N5578, N5514, N5515);
nor NOR2_2095 (N5581, N5519, N5516);
nor NOR2_2096 (N5585, N5464, N5522);
nor NOR2_2097 (N5586, N5522, N5461);
nor NOR2_2098 (N5587, N5526, N5527);
nor NOR2_2099 (N5590, N5528, N1164);
nor NOR2_2100 (N5594, N5473, N5531);
nor NOR2_2101 (N5595, N5531, N1212);
nor NOR2_2102 (N5596, N5360, N5531);
nor NOR2_2103 (N5599, N5535, N5536);
nor NOR2_2104 (N5602, N1308, N5537);
nor NOR2_2105 (N5606, N5480, N5540);
nor NOR2_2106 (N5607, N5540, N582);
nor NOR2_2107 (N5608, N5366, N5540);
nor NOR2_2108 (N5611, N5483, N5544);
nor NOR2_2109 (N5612, N5544, N630);
nor NOR2_2110 (N5613, N5370, N5544);
nor NOR2_2111 (N5616, N5486, N5548);
nor NOR2_2112 (N5617, N5548, N678);
nor NOR2_2113 (N5618, N5374, N5548);
nor NOR2_2114 (N5621, N5552, N5553);
  nor NOR2_2115 (keyinput_Wire_0[252], N5557, N5554);
  xor keyGate_0_252(KeyNOTWire_0[139], keyinput252, keyinput_Wire_0[252]);
  not KeyNOTGate_0_139(N5624, KeyNOTWire_0[139]);
nor NOR2_2116 (N5628, N5498, N5560);
nor NOR2_2117 (N5629, N5560, N5495);
nor NOR2_2118 (N5630, N5564, N5565);
nor NOR2_2119 (N5633, N5566, N873);
nor NOR2_2120 (N5637, N5507, N5569);
nor NOR2_2121 (N5638, N5569, N921);
nor NOR2_2122 (N5639, N5395, N5569);
nor NOR2_2123 (N5642, N5573, N5574);
nor NOR2_2124 (N5645, N5578, N5575);
nor NOR2_2125 (N5649, N5519, N5581);
nor NOR2_2126 (N5650, N5581, N5516);
nor NOR2_2127 (N5651, N5585, N5586);
nor NOR2_2128 (N5654, N5587, N1116);
nor NOR2_2129 (N5658, N5528, N5590);
nor NOR2_2130 (N5659, N5590, N1164);
nor NOR2_2131 (N5660, N5416, N5590);
nor NOR2_2132 (N5663, N5594, N5595);
nor NOR2_2133 (N5666, N5599, N5596);
nor NOR2_2134 (N5670, N1308, N5602);
nor NOR2_2135 (N5671, N5602, N5537);
nor NOR2_2136 (N5672, N5606, N5607);
nor NOR2_2137 (N5673, N5611, N5612);
nor NOR2_2138 (N5676, N5616, N5617);
nor NOR2_2139 (N5679, N5621, N5618);
nor NOR2_2140 (N5683, N5557, N5624);
nor NOR2_2141 (N5684, N5624, N5554);
nor NOR2_2142 (N5685, N5628, N5629);
nor NOR2_2143 (N5688, N5630, N825);
nor NOR2_2144 (N5692, N5566, N5633);
nor NOR2_2145 (N5693, N5633, N873);
nor NOR2_2146 (N5694, N5446, N5633);
nor NOR2_2147 (N5697, N5637, N5638);
nor NOR2_2148 (N5700, N5642, N5639);
nor NOR2_2149 (N5704, N5578, N5645);
nor NOR2_2150 (N5705, N5645, N5575);
nor NOR2_2151 (N5706, N5649, N5650);
nor NOR2_2152 (N5709, N5651, N1068);
nor NOR2_2153 (N5713, N5587, N5654);
nor NOR2_2154 (N5714, N5654, N1116);
nor NOR2_2155 (N5715, N5467, N5654);
nor NOR2_2156 (N5718, N5658, N5659);
nor NOR2_2157 (N5721, N5663, N5660);
nor NOR2_2158 (N5725, N5599, N5666);
nor NOR2_2159 (N5726, N5666, N5596);
nor NOR2_2160 (N5727, N5670, N5671);
nor NOR2_2161 (N5730, N5673, N5608);
nor NOR2_2162 (N5734, N5676, N5613);
nor NOR2_2163 (N5738, N5621, N5679);
nor NOR2_2164 (N5739, N5679, N5618);
nor NOR2_2165 (N5740, N5683, N5684);
nor NOR2_2166 (N5743, N5685, N777);
nor NOR2_2167 (N5747, N5630, N5688);
nor NOR2_2168 (N5748, N5688, N825);
nor NOR2_2169 (N5749, N5501, N5688);
nor NOR2_2170 (N5752, N5692, N5693);
nor NOR2_2171 (N5755, N5697, N5694);
nor NOR2_2172 (N5759, N5642, N5700);
nor NOR2_2173 (N5760, N5700, N5639);
nor NOR2_2174 (N5761, N5704, N5705);
nor NOR2_2175 (N5764, N5706, N1020);
nor NOR2_2176 (N5768, N5651, N5709);
nor NOR2_2177 (N5769, N5709, N1068);
nor NOR2_2178 (N5770, N5522, N5709);
nor NOR2_2179 (N5773, N5713, N5714);
nor NOR2_2180 (N5776, N5718, N5715);
nor NOR2_2181 (N5780, N5663, N5721);
nor NOR2_2182 (N5781, N5721, N5660);
nor NOR2_2183 (N5782, N5725, N5726);
nor NOR2_2184 (N5785, N5673, N5730);
nor NOR2_2185 (N5786, N5730, N5608);
nor NOR2_2186 (N5787, N5676, N5734);
nor NOR2_2187 (N5788, N5734, N5613);
nor NOR2_2188 (N5789, N5738, N5739);
nor NOR2_2189 (N5792, N5740, N729);
nor NOR2_2190 (N5796, N5685, N5743);
nor NOR2_2191 (N5797, N5743, N777);
nor NOR2_2192 (N5798, N5560, N5743);
nor NOR2_2193 (N5801, N5747, N5748);
nor NOR2_2194 (N5804, N5752, N5749);
nor NOR2_2195 (N5808, N5697, N5755);
nor NOR2_2196 (N5809, N5755, N5694);
nor NOR2_2197 (N5810, N5759, N5760);
nor NOR2_2198 (N5813, N5761, N972);
nor NOR2_2199 (N5817, N5706, N5764);
nor NOR2_2200 (N5818, N5764, N1020);
nor NOR2_2201 (N5819, N5581, N5764);
nor NOR2_2202 (N5822, N5768, N5769);
nor NOR2_2203 (N5825, N5773, N5770);
nor NOR2_2204 (N5829, N5718, N5776);
nor NOR2_2205 (N5830, N5776, N5715);
nor NOR2_2206 (N5831, N5780, N5781);
nor NOR2_2207 (N5834, N5785, N5786);
nor NOR2_2208 (N5837, N5787, N5788);
nor NOR2_2209 (N5840, N5789, N681);
nor NOR2_2210 (N5844, N5740, N5792);
nor NOR2_2211 (N5845, N5792, N729);
nor NOR2_2212 (N5846, N5624, N5792);
nor NOR2_2213 (N5849, N5796, N5797);
nor NOR2_2214 (N5852, N5801, N5798);
nor NOR2_2215 (N5856, N5752, N5804);
nor NOR2_2216 (N5857, N5804, N5749);
nor NOR2_2217 (N5858, N5808, N5809);
nor NOR2_2218 (N5861, N5810, N924);
nor NOR2_2219 (N5865, N5761, N5813);
nor NOR2_2220 (N5866, N5813, N972);
nor NOR2_2221 (N5867, N5645, N5813);
nor NOR2_2222 (N5870, N5817, N5818);
nor NOR2_2223 (N5873, N5822, N5819);
nor NOR2_2224 (N5877, N5773, N5825);
nor NOR2_2225 (N5878, N5825, N5770);
nor NOR2_2226 (N5879, N5829, N5830);
nor NOR2_2227 (N5882, N5834, N585);
nor NOR2_2228 (N5886, N5837, N633);
nor NOR2_2229 (N5890, N5789, N5840);
nor NOR2_2230 (N5891, N5840, N681);
nor NOR2_2231 (N5892, N5679, N5840);
nor NOR2_2232 (N5895, N5844, N5845);
nor NOR2_2233 (N5898, N5849, N5846);
nor NOR2_2234 (N5902, N5801, N5852);
nor NOR2_2235 (N5903, N5852, N5798);
nor NOR2_2236 (N5904, N5856, N5857);
nor NOR2_2237 (N5907, N5858, N876);
nor NOR2_2238 (N5911, N5810, N5861);
  nor NOR2_2239 (keyinput_Wire_0[253], N5861, N924);
  xnor keyGate_0_253(KeyNOTWire_0[140], keyinput253, keyinput_Wire_0[253]);
  not KeyNOTGate_0_140(N5912, KeyNOTWire_0[140]);
nor NOR2_2240 (N5913, N5700, N5861);
nor NOR2_2241 (N5916, N5865, N5866);
nor NOR2_2242 (N5919, N5870, N5867);
nor NOR2_2243 (N5923, N5822, N5873);
nor NOR2_2244 (N5924, N5873, N5819);
nor NOR2_2245 (N5925, N5877, N5878);
nor NOR2_2246 (N5928, N5834, N5882);
nor NOR2_2247 (N5929, N5882, N585);
nor NOR2_2248 (N5930, N5730, N5882);
nor NOR2_2249 (N5933, N5837, N5886);
nor NOR2_2250 (N5934, N5886, N633);
nor NOR2_2251 (N5935, N5734, N5886);
nor NOR2_2252 (N5938, N5890, N5891);
nor NOR2_2253 (N5941, N5895, N5892);
nor NOR2_2254 (N5945, N5849, N5898);
nor NOR2_2255 (N5946, N5898, N5846);
nor NOR2_2256 (N5947, N5902, N5903);
nor NOR2_2257 (N5950, N5904, N828);
nor NOR2_2258 (N5954, N5858, N5907);
nor NOR2_2259 (N5955, N5907, N876);
nor NOR2_2260 (N5956, N5755, N5907);
nor NOR2_2261 (N5959, N5911, N5912);
nor NOR2_2262 (N5962, N5916, N5913);
nor NOR2_2263 (N5966, N5870, N5919);
nor NOR2_2264 (N5967, N5919, N5867);
nor NOR2_2265 (N5968, N5923, N5924);
nor NOR2_2266 (N5971, N5928, N5929);
nor NOR2_2267 (N5972, N5933, N5934);
nor NOR2_2268 (N5975, N5938, N5935);
nor NOR2_2269 (N5979, N5895, N5941);
nor NOR2_2270 (N5980, N5941, N5892);
nor NOR2_2271 (N5981, N5945, N5946);
nor NOR2_2272 (N5984, N5947, N780);
nor NOR2_2273 (N5988, N5904, N5950);
nor NOR2_2274 (N5989, N5950, N828);
nor NOR2_2275 (N5990, N5804, N5950);
nor NOR2_2276 (N5993, N5954, N5955);
nor NOR2_2277 (N5996, N5959, N5956);
nor NOR2_2278 (N6000, N5916, N5962);
nor NOR2_2279 (N6001, N5962, N5913);
nor NOR2_2280 (N6002, N5966, N5967);
nor NOR2_2281 (N6005, N5972, N5930);
nor NOR2_2282 (N6009, N5938, N5975);
nor NOR2_2283 (N6010, N5975, N5935);
nor NOR2_2284 (N6011, N5979, N5980);
nor NOR2_2285 (N6014, N5981, N732);
nor NOR2_2286 (N6018, N5947, N5984);
nor NOR2_2287 (N6019, N5984, N780);
nor NOR2_2288 (N6020, N5852, N5984);
nor NOR2_2289 (N6023, N5988, N5989);
nor NOR2_2290 (N6026, N5993, N5990);
nor NOR2_2291 (N6030, N5959, N5996);
nor NOR2_2292 (N6031, N5996, N5956);
nor NOR2_2293 (N6032, N6000, N6001);
nor NOR2_2294 (N6035, N5972, N6005);
nor NOR2_2295 (N6036, N6005, N5930);
nor NOR2_2296 (N6037, N6009, N6010);
nor NOR2_2297 (N6040, N6011, N684);
nor NOR2_2298 (N6044, N5981, N6014);
nor NOR2_2299 (N6045, N6014, N732);
nor NOR2_2300 (N6046, N5898, N6014);
nor NOR2_2301 (N6049, N6018, N6019);
nor NOR2_2302 (N6052, N6023, N6020);
nor NOR2_2303 (N6056, N5993, N6026);
nor NOR2_2304 (N6057, N6026, N5990);
nor NOR2_2305 (N6058, N6030, N6031);
nor NOR2_2306 (N6061, N6035, N6036);
nor NOR2_2307 (N6064, N6037, N636);
nor NOR2_2308 (N6068, N6011, N6040);
nor NOR2_2309 (N6069, N6040, N684);
nor NOR2_2310 (N6070, N5941, N6040);
nor NOR2_2311 (N6073, N6044, N6045);
nor NOR2_2312 (N6076, N6049, N6046);
nor NOR2_2313 (N6080, N6023, N6052);
nor NOR2_2314 (N6081, N6052, N6020);
nor NOR2_2315 (N6082, N6056, N6057);
nor NOR2_2316 (N6085, N6061, N588);
nor NOR2_2317 (N6089, N6037, N6064);
nor NOR2_2318 (N6090, N6064, N636);
nor NOR2_2319 (N6091, N5975, N6064);
nor NOR2_2320 (N6094, N6068, N6069);
nor NOR2_2321 (N6097, N6073, N6070);
nor NOR2_2322 (N6101, N6049, N6076);
nor NOR2_2323 (N6102, N6076, N6046);
nor NOR2_2324 (N6103, N6080, N6081);
nor NOR2_2325 (N6106, N6061, N6085);
nor NOR2_2326 (N6107, N6085, N588);
nor NOR2_2327 (N6108, N6005, N6085);
nor NOR2_2328 (N6111, N6089, N6090);
nor NOR2_2329 (N6114, N6094, N6091);
nor NOR2_2330 (N6118, N6073, N6097);
nor NOR2_2331 (N6119, N6097, N6070);
nor NOR2_2332 (N6120, N6101, N6102);
nor NOR2_2333 (N6123, N6106, N6107);
  nor NOR2_2334 (keyinput_Wire_0[254], N6111, N6108);
  xor keyGate_0_254(KeyNOTWire_0[141], keyinput254, keyinput_Wire_0[254]);
  not KeyNOTGate_0_141(N6124, KeyNOTWire_0[141]);
nor NOR2_2335 (N6128, N6094, N6114);
nor NOR2_2336 (N6129, N6114, N6091);
nor NOR2_2337 (N6130, N6118, N6119);
nor NOR2_2338 (N6133, N6111, N6124);
nor NOR2_2339 (N6134, N6124, N6108);
nor NOR2_2340 (N6135, N6128, N6129);
nor NOR2_2341 (N6138, N6133, N6134);
not NOT1_2342 (N6141, N6138);
nor NOR2_2343 (N6145, N6138, N6141);
not NOT1_2344 (N6146, N6141);
nor NOR2_2345 (N6147, N6124, N6141);
nor NOR2_2346 (N6150, N6145, N6146);
nor NOR2_2347 (N6151, N6135, N6147);
nor NOR2_2348 (N6155, N6135, N6151);
nor NOR2_2349 (N6156, N6151, N6147);
nor NOR2_2350 (N6157, N6114, N6151);
nor NOR2_2351 (N6160, N6155, N6156);
nor NOR2_2352 (N6161, N6130, N6157);
nor NOR2_2353 (N6165, N6130, N6161);
nor NOR2_2354 (N6166, N6161, N6157);
nor NOR2_2355 (N6167, N6097, N6161);
nor NOR2_2356 (N6170, N6165, N6166);
nor NOR2_2357 (N6171, N6120, N6167);
nor NOR2_2358 (N6175, N6120, N6171);
nor NOR2_2359 (N6176, N6171, N6167);
nor NOR2_2360 (N6177, N6076, N6171);
nor NOR2_2361 (N6180, N6175, N6176);
nor NOR2_2362 (N6181, N6103, N6177);
nor NOR2_2363 (N6185, N6103, N6181);
nor NOR2_2364 (N6186, N6181, N6177);
nor NOR2_2365 (N6187, N6052, N6181);
nor NOR2_2366 (N6190, N6185, N6186);
nor NOR2_2367 (N6191, N6082, N6187);
nor NOR2_2368 (N6195, N6082, N6191);
nor NOR2_2369 (N6196, N6191, N6187);
nor NOR2_2370 (N6197, N6026, N6191);
nor NOR2_2371 (N6200, N6195, N6196);
nor NOR2_2372 (N6201, N6058, N6197);
nor NOR2_2373 (N6205, N6058, N6201);
nor NOR2_2374 (N6206, N6201, N6197);
nor NOR2_2375 (N6207, N5996, N6201);
  nor NOR2_2376 (keyinput_Wire_0[255], N6205, N6206);
  xnor keyGate_0_255(KeyNOTWire_0[142], keyinput255, keyinput_Wire_0[255]);
  not KeyNOTGate_0_142(N6210, KeyNOTWire_0[142]);
nor NOR2_2377 (N6211, N6032, N6207);
nor NOR2_2378 (N6215, N6032, N6211);
nor NOR2_2379 (N6216, N6211, N6207);
nor NOR2_2380 (N6217, N5962, N6211);
nor NOR2_2381 (N6220, N6215, N6216);
nor NOR2_2382 (N6221, N6002, N6217);
nor NOR2_2383 (N6225, N6002, N6221);
nor NOR2_2384 (N6226, N6221, N6217);
nor NOR2_2385 (N6227, N5919, N6221);
nor NOR2_2386 (N6230, N6225, N6226);
nor NOR2_2387 (N6231, N5968, N6227);
nor NOR2_2388 (N6235, N5968, N6231);
nor NOR2_2389 (N6236, N6231, N6227);
nor NOR2_2390 (N6237, N5873, N6231);
nor NOR2_2391 (N6240, N6235, N6236);
nor NOR2_2392 (N6241, N5925, N6237);
nor NOR2_2393 (N6245, N5925, N6241);
nor NOR2_2394 (N6246, N6241, N6237);
nor NOR2_2395 (N6247, N5825, N6241);
nor NOR2_2396 (N6250, N6245, N6246);
nor NOR2_2397 (N6251, N5879, N6247);
nor NOR2_2398 (N6255, N5879, N6251);
nor NOR2_2399 (N6256, N6251, N6247);
nor NOR2_2400 (N6257, N5776, N6251);
nor NOR2_2401 (N6260, N6255, N6256);
nor NOR2_2402 (N6261, N5831, N6257);
nor NOR2_2403 (N6265, N5831, N6261);
nor NOR2_2404 (N6266, N6261, N6257);
nor NOR2_2405 (N6267, N5721, N6261);
nor NOR2_2406 (N6270, N6265, N6266);
nor NOR2_2407 (N6271, N5782, N6267);
nor NOR2_2408 (N6275, N5782, N6271);
nor NOR2_2409 (N6276, N6271, N6267);
nor NOR2_2410 (N6277, N5666, N6271);
nor NOR2_2411 (N6280, N6275, N6276);
nor NOR2_2412 (N6281, N5727, N6277);
nor NOR2_2413 (N6285, N5727, N6281);
nor NOR2_2414 (N6286, N6281, N6277);
nor NOR2_2415 (N6287, N5602, N6281);
nor NOR2_2416 (N6288, N6285, N6286);

AntiSAT some_name( KeyWire_0_2, N341, N1, N528, N443, N375, N307, N120, N171, N52, N426, N18, N460, N256, N154, N324, N290, N494, N239, N477, N392, N137, N103, N86, N205, N273, N69, N409, N511, N222, N188, N358, N35, keyinput256, keyinput257, keyinput258, keyinput259, keyinput260, keyinput261, keyinput262, keyinput263, keyinput264, keyinput265, keyinput266, keyinput267, keyinput268, keyinput269, keyinput270, keyinput271, keyinput272, keyinput273, keyinput274, keyinput275, keyinput276, keyinput277, keyinput278, keyinput279, keyinput280, keyinput281, keyinput282, keyinput283, keyinput284, keyinput285, keyinput286, keyinput287, keyinput288, keyinput289, keyinput290, keyinput291, keyinput292, keyinput293, keyinput294, keyinput295, keyinput296, keyinput297, keyinput298, keyinput299, keyinput300, keyinput301, keyinput302, keyinput303, keyinput304, keyinput305, keyinput306, keyinput307, keyinput308, keyinput309, keyinput310, keyinput311, keyinput312, keyinput313, keyinput314, keyinput315, keyinput316, keyinput317, keyinput318, keyinput319,
       keyinput320, keyinput321, keyinput322, keyinput323, keyinput324,
       keyinput325, keyinput326, keyinput327, keyinput328, keyinput329,
       keyinput330, keyinput331, keyinput332, keyinput333, keyinput334,
       keyinput335, keyinput336, keyinput337, keyinput338, keyinput339,
       keyinput340, keyinput341, keyinput342, keyinput343, keyinput344,
       keyinput345, keyinput346, keyinput347, keyinput348, keyinput349,
       keyinput350, keyinput351);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N341, N1, N528, N443, N375, N307, N120, N171, N52, N426, N18, N460, N256, N154, N324, N290, N494, N239, N477, N392, N137, N103, N86, N205, N273, N69, N409, N511, N222, N188, N358, N35, keyinput256, keyinput257, keyinput258, keyinput259, keyinput260, keyinput261, keyinput262, keyinput263, keyinput264, keyinput265, keyinput266, keyinput267, keyinput268, keyinput269, keyinput270, keyinput271, keyinput272, keyinput273, keyinput274, keyinput275, keyinput276, keyinput277, keyinput278, keyinput279, keyinput280, keyinput281, keyinput282, keyinput283, keyinput284, keyinput285, keyinput286, keyinput287, keyinput288, keyinput289, keyinput290, keyinput291, keyinput292, keyinput293, keyinput294, keyinput295, keyinput296, keyinput297, keyinput298, keyinput299, keyinput300, keyinput301, keyinput302, keyinput303, keyinput304, keyinput305, keyinput306, keyinput307, keyinput308, keyinput309, keyinput310, keyinput311, keyinput312, keyinput313, keyinput314, keyinput315, keyinput316, keyinput317, keyinput318, keyinput319 ,
        keyinput320, keyinput321, keyinput322, keyinput323, keyinput324,
        keyinput325, keyinput326, keyinput327, keyinput328, keyinput329,
        keyinput330, keyinput331, keyinput332, keyinput333, keyinput334,
        keyinput335, keyinput336, keyinput337, keyinput338, keyinput339,
        keyinput340, keyinput341, keyinput342, keyinput343, keyinput344,
        keyinput345, keyinput346, keyinput347, keyinput348, keyinput349,
        keyinput350, keyinput351);

  input keyinput320, keyinput321, keyinput322, keyinput323, keyinput324;
  input keyinput325, keyinput326, keyinput327, keyinput328, keyinput329;
  input keyinput330, keyinput331, keyinput332, keyinput333, keyinput334;
  input keyinput335, keyinput336, keyinput337, keyinput338, keyinput339;
  input keyinput340, keyinput341, keyinput342, keyinput343, keyinput344;
  input keyinput345, keyinput346, keyinput347, keyinput348, keyinput349;
  input keyinput350, keyinput351;

  wire [0:31] keyNTin_Wire_1;
  wire [0:18] KeyNOTWire_1;

  input N341, N1, N528, N443, N375, N307, N120, N171, N52, N426, N18, N460, N256, N154, N324, N290, N494, N239, N477, N392, N137, N103, N86, N205, N273, N69, N409, N511, N222, N188, N358, N35;
  input keyinput256, keyinput257, keyinput258, keyinput259, keyinput260, keyinput261, keyinput262, keyinput263, keyinput264, keyinput265, keyinput266, keyinput267, keyinput268, keyinput269, keyinput270, keyinput271, keyinput272, keyinput273, keyinput274, keyinput275, keyinput276, keyinput277, keyinput278, keyinput279, keyinput280, keyinput281, keyinput282, keyinput283, keyinput284, keyinput285, keyinput286, keyinput287, keyinput288, keyinput289, keyinput290, keyinput291, keyinput292, keyinput293, keyinput294, keyinput295, keyinput296, keyinput297, keyinput298, keyinput299, keyinput300, keyinput301, keyinput302, keyinput303, keyinput304, keyinput305, keyinput306, keyinput307, keyinput308, keyinput309, keyinput310, keyinput311, keyinput312, keyinput313, keyinput314, keyinput315, keyinput316, keyinput317, keyinput318, keyinput319;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65 ;

  xnor KeyGate0 (keyNTin_Wire_1[0], N341, keyinput256);
  xor keyNTinGate_1_0(KeyNOTWire_1[0], keyinput320, keyNTin_Wire_1[0]);
  not KeyNOTGate_1_0(newWire_0, KeyNOTWire_1[0]);
  xor  KeyGate1 (newWire_1, N1, keyinput257);
  xnor KeyGate2 (keyNTin_Wire_1[1], N528, keyinput258);
  xor keyNTinGate_1_1(KeyNOTWire_1[1], keyinput321, keyNTin_Wire_1[1]);
  not KeyNOTGate_1_1(newWire_2, KeyNOTWire_1[1]);
  xnor KeyGate3 (newWire_3, N443, keyinput259);
  xor  KeyGate4 (keyNTin_Wire_1[2], N375, keyinput260);
  xor keyNTinGate_1_2(newWire_4, keyinput322, keyNTin_Wire_1[2]);
  xor  KeyGate5 (keyNTin_Wire_1[3], N307, keyinput261);
  xor keyNTinGate_1_3(newWire_5, keyinput323, keyNTin_Wire_1[3]);
  xor  KeyGate6 (newWire_6, N120, keyinput262);
  xor  KeyGate7 (newWire_7, N171, keyinput263);
  xnor KeyGate8 (newWire_8, N52, keyinput264);
  xor  KeyGate9 (keyNTin_Wire_1[4], N426, keyinput265);
  xnor keyNTinGate_1_4(KeyNOTWire_1[2], keyinput324, keyNTin_Wire_1[4]);
  not KeyNOTGate_1_2(newWire_9, KeyNOTWire_1[2]);
  xor  KeyGate10 (keyNTin_Wire_1[5], N18, keyinput266);
  xor keyNTinGate_1_5(newWire_10, keyinput325, keyNTin_Wire_1[5]);
  xnor KeyGate11 (keyNTin_Wire_1[6], N460, keyinput267);
  xor keyNTinGate_1_6(newWire_11, keyinput326, keyNTin_Wire_1[6]);
  xor  KeyGate12 (keyNTin_Wire_1[7], N256, keyinput268);
  xor keyNTinGate_1_7(KeyNOTWire_1[3], keyinput327, keyNTin_Wire_1[7]);
  not KeyNOTGate_1_3(newWire_12, KeyNOTWire_1[3]);
  xor  KeyGate13 (newWire_13, N154, keyinput269);
  xor  KeyGate14 (newWire_14, N324, keyinput270);
  xnor KeyGate15 (newWire_15, N290, keyinput271);
  xor  KeyGate16 (keyNTin_Wire_1[8], N494, keyinput272);
  xor keyNTinGate_1_8(KeyNOTWire_1[4], keyinput328, keyNTin_Wire_1[8]);
  not KeyNOTGate_1_4(newWire_16, KeyNOTWire_1[4]);
  xnor KeyGate17 (keyNTin_Wire_1[9], N239, keyinput273);
  xnor keyNTinGate_1_9(KeyNOTWire_1[5], keyinput329, keyNTin_Wire_1[9]);
  not KeyNOTGate_1_5(newWire_17, KeyNOTWire_1[5]);
  xor  KeyGate18 (keyNTin_Wire_1[10], N477, keyinput274);
  xnor keyNTinGate_1_10(KeyNOTWire_1[6], keyinput330, keyNTin_Wire_1[10]);
  not KeyNOTGate_1_6(newWire_18, KeyNOTWire_1[6]);
  xnor KeyGate19 (newWire_19, N392, keyinput275);
  xnor KeyGate20 (keyNTin_Wire_1[11], N137, keyinput276);
  xor keyNTinGate_1_11(KeyNOTWire_1[7], keyinput331, keyNTin_Wire_1[11]);
  not KeyNOTGate_1_7(newWire_20, KeyNOTWire_1[7]);
  xnor KeyGate21 (newWire_21, N103, keyinput277);
  xor  KeyGate22 (newWire_22, N86, keyinput278);
  xor  KeyGate23 (keyNTin_Wire_1[12], N205, keyinput279);
  xnor keyNTinGate_1_12(KeyNOTWire_1[8], keyinput332, keyNTin_Wire_1[12]);
  not KeyNOTGate_1_8(newWire_23, KeyNOTWire_1[8]);
  xnor KeyGate24 (newWire_24, N273, keyinput280);
  xor  KeyGate25 (newWire_25, N69, keyinput281);
  xnor KeyGate26 (newWire_26, N409, keyinput282);
  xor  KeyGate27 (newWire_27, N511, keyinput283);
  xnor KeyGate28 (newWire_28, N222, keyinput284);
  xnor KeyGate29 (keyNTin_Wire_1[13], N188, keyinput285);
  xnor keyNTinGate_1_13(newWire_29, keyinput333, keyNTin_Wire_1[13]);
  xor  KeyGate30 (keyNTin_Wire_1[14], N358, keyinput286);
  xnor keyNTinGate_1_14(KeyNOTWire_1[9], keyinput334, keyNTin_Wire_1[14]);
  not KeyNOTGate_1_9(newWire_30, KeyNOTWire_1[9]);
  xnor KeyGate31 (keyNTin_Wire_1[15], N35, keyinput287);
  xnor keyNTinGate_1_15(KeyNOTWire_1[10], keyinput335, keyNTin_Wire_1[15]);
  not KeyNOTGate_1_10(newWire_31, KeyNOTWire_1[10]);
  xnor KeyGate32 (newWire_32, N341, keyinput288);
  xnor KeyGate33 (newWire_33, N1, keyinput289);
  xnor KeyGate34 (keyNTin_Wire_1[16], N528, keyinput290);
  xor keyNTinGate_1_16(newWire_34, keyinput336, keyNTin_Wire_1[16]);
  xnor KeyGate35 (newWire_35, N443, keyinput291);
  xor  KeyGate36 (keyNTin_Wire_1[17], N375, keyinput292);
  xor keyNTinGate_1_17(KeyNOTWire_1[11], keyinput337, keyNTin_Wire_1[17]);
  not KeyNOTGate_1_11(newWire_36, KeyNOTWire_1[11]);
  xnor KeyGate37 (newWire_37, N307, keyinput293);
  xnor KeyGate38 (newWire_38, N120, keyinput294);
  xnor KeyGate39 (newWire_39, N171, keyinput295);
  xor  KeyGate40 (newWire_40, N52, keyinput296);
  xnor KeyGate41 (keyNTin_Wire_1[18], N426, keyinput297);
  xor keyNTinGate_1_18(KeyNOTWire_1[12], keyinput338, keyNTin_Wire_1[18]);
  not KeyNOTGate_1_12(newWire_41, KeyNOTWire_1[12]);
  xor  KeyGate42 (newWire_42, N18, keyinput298);
  xor  KeyGate43 (keyNTin_Wire_1[19], N460, keyinput299);
  xor keyNTinGate_1_19(newWire_43, keyinput339, keyNTin_Wire_1[19]);
  xor  KeyGate44 (keyNTin_Wire_1[20], N256, keyinput300);
  xor keyNTinGate_1_20(newWire_44, keyinput340, keyNTin_Wire_1[20]);
  xnor KeyGate45 (keyNTin_Wire_1[21], N154, keyinput301);
  xor keyNTinGate_1_21(KeyNOTWire_1[13], keyinput341, keyNTin_Wire_1[21]);
  not KeyNOTGate_1_13(newWire_45, KeyNOTWire_1[13]);
  xnor KeyGate46 (keyNTin_Wire_1[22], N324, keyinput302);
  xor keyNTinGate_1_22(newWire_46, keyinput342, keyNTin_Wire_1[22]);
  xnor KeyGate47 (keyNTin_Wire_1[23], N290, keyinput303);
  xnor keyNTinGate_1_23(KeyNOTWire_1[14], keyinput343, keyNTin_Wire_1[23]);
  not KeyNOTGate_1_14(newWire_47, KeyNOTWire_1[14]);
  xnor KeyGate48 (keyNTin_Wire_1[24], N494, keyinput304);
  xor keyNTinGate_1_24(newWire_48, keyinput344, keyNTin_Wire_1[24]);
  xnor KeyGate49 (keyNTin_Wire_1[25], N239, keyinput305);
  xor keyNTinGate_1_25(KeyNOTWire_1[15], keyinput345, keyNTin_Wire_1[25]);
  not KeyNOTGate_1_15(newWire_49, KeyNOTWire_1[15]);
  xor  KeyGate50 (keyNTin_Wire_1[26], N477, keyinput306);
  xor keyNTinGate_1_26(newWire_50, keyinput346, keyNTin_Wire_1[26]);
  xor  KeyGate51 (newWire_51, N392, keyinput307);
  xnor KeyGate52 (keyNTin_Wire_1[27], N137, keyinput308);
  xor keyNTinGate_1_27(newWire_52, keyinput347, keyNTin_Wire_1[27]);
  xnor KeyGate53 (keyNTin_Wire_1[28], N103, keyinput309);
  xor keyNTinGate_1_28(newWire_53, keyinput348, keyNTin_Wire_1[28]);
  xnor KeyGate54 (newWire_54, N86, keyinput310);
  xor  KeyGate55 (newWire_55, N205, keyinput311);
  xor  KeyGate56 (keyNTin_Wire_1[29], N273, keyinput312);
  xor keyNTinGate_1_29(KeyNOTWire_1[16], keyinput349, keyNTin_Wire_1[29]);
  not KeyNOTGate_1_16(newWire_56, KeyNOTWire_1[16]);
  xnor KeyGate57 (newWire_57, N69, keyinput313);
  xnor KeyGate58 (keyNTin_Wire_1[30], N409, keyinput314);
  xnor keyNTinGate_1_30(KeyNOTWire_1[17], keyinput350, keyNTin_Wire_1[30]);
  not KeyNOTGate_1_17(newWire_58, KeyNOTWire_1[17]);
  xnor KeyGate59 (newWire_59, N511, keyinput315);
  xor  KeyGate60 (newWire_60, N222, keyinput316);
  xnor KeyGate61 (newWire_61, N188, keyinput317);
  xnor KeyGate62 (newWire_62, N358, keyinput318);
  xnor KeyGate63 (newWire_63, N35, keyinput319);
  and some_function (keyNTin_Wire_1[31], newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31 );
  xor keyNTinGate_1_31(KeyNOTWire_1[18], keyinput351, keyNTin_Wire_1[31]);
  not KeyNOTGate_1_18(newWire_64, KeyNOTWire_1[18]);
  nand compl_function (newWire_65, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63);
  and finalAND (KeyWire_0_2, newWire_64, newWire_65);

endmodule /* AntiSAT */
