// Verilog File 
module top (G1gat,G8gat,G13gat,G17gat,G26gat,G29gat,G36gat,G42gat,G51gat,
G55gat,G59gat,G68gat,G72gat,G73gat,G74gat,G75gat,G80gat,G85gat,G86gat,
G87gat,G88gat,G89gat,G90gat,G91gat,G96gat,G101gat,G106gat,G111gat,G116gat,
G121gat,G126gat,G130gat,G135gat,G138gat,G143gat,G146gat,G149gat,G152gat,G153gat,
G156gat,G159gat,G165gat,G171gat,G177gat,G183gat,G189gat,G195gat,G201gat,G207gat,
G210gat,G219gat,G228gat,G237gat,G246gat,G255gat,G259gat,G260gat,G261gat,G267gat,
G268gat,G388gat,G389gat,G390gat,G391gat,G418gat,G419gat,G420gat,G421gat,G422gat,
G423gat,G446gat,G447gat,G448gat,G449gat,G450gat,G767gat,G768gat,G850gat,G863gat,
G864gat,G865gat,G866gat,G874gat,G878gat,G879gat,G880gat,keyinput0,keyinput1,keyinput2,
keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,
keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,
keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,
keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,
keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,
keyinput53,keyinput54,keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,
keyinput63,keyinput64,keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,
keyinput73,keyinput74,keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,
keyinput83,keyinput84,keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,
keyinput93,keyinput94,keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,
keyinput103,keyinput104,keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,
keyinput113,keyinput114,keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,
keyinput123,keyinput124,keyinput125,keyinput126,keyinput127,keyinput128,keyinput129,keyinput130,keyinput131,keyinput132,
keyinput133,keyinput134,keyinput135,keyinput136,keyinput137,keyinput138,keyinput139,keyinput140,keyinput141,keyinput142,
keyinput143,keyinput144,keyinput145,keyinput146,keyinput147,keyinput148,keyinput149,keyinput150,keyinput151,keyinput152,
keyinput153,keyinput154,keyinput155,keyinput156,keyinput157,keyinput158,keyinput159,keyinput160,keyinput161,keyinput162,
keyinput163,keyinput164,keyinput165,keyinput166,keyinput167,keyinput168,keyinput169,keyinput170,keyinput171,keyinput172,
keyinput173,keyinput174,keyinput175,keyinput176,keyinput177,keyinput178,keyinput179,keyinput180,keyinput181,keyinput182,
keyinput183,keyinput184,keyinput185,keyinput186,keyinput187,keyinput188,keyinput189,keyinput190,keyinput191,keyinput192,
keyinput193,keyinput194,keyinput195,keyinput196,keyinput197,keyinput198,keyinput199,keyinput200,keyinput201,keyinput202,
keyinput203,keyinput204,keyinput205,keyinput206,keyinput207,keyinput208,keyinput209,keyinput210,keyinput211,keyinput212,
keyinput213,keyinput214,keyinput215,keyinput216,keyinput217,keyinput218,keyinput219,keyinput220,keyinput221,keyinput222,
keyinput223,keyinput224,keyinput225,keyinput226,keyinput227,keyinput228,keyinput229,keyinput230,keyinput231,keyinput232,
keyinput233,keyinput234,keyinput235,keyinput236,keyinput237,keyinput238,keyinput239,keyinput240,keyinput241,keyinput242,
keyinput243,keyinput244,keyinput245,keyinput246,keyinput247,keyinput248,keyinput249,keyinput250,keyinput251,keyinput252,
keyinput253,keyinput254,keyinput255,keyinput256,keyinput257,keyinput258,keyinput259,keyinput260,keyinput261,keyinput262,
keyinput263,keyinput264,keyinput265,keyinput266,keyinput267,keyinput268,keyinput269,keyinput270,keyinput271,keyinput272,
keyinput273,keyinput274,keyinput275,keyinput276,keyinput277,keyinput278,keyinput279,keyinput280,keyinput281,keyinput282,
keyinput283,keyinput284,keyinput285,keyinput286,keyinput287,keyinput288,keyinput289,keyinput290,keyinput291,keyinput292,
keyinput293,keyinput294,keyinput295,keyinput296,keyinput297,keyinput298,keyinput299,keyinput300,keyinput301,keyinput302,
keyinput303,keyinput304,keyinput305,keyinput306,keyinput307,keyinput308,keyinput309,keyinput310,keyinput311,keyinput312,
keyinput313,keyinput314,keyinput315,keyinput316,keyinput317,keyinput318,keyinput319,keyinput320,keyinput321,keyinput322,
keyinput323,keyinput324,keyinput325,keyinput326,keyinput327,keyinput328,keyinput329,keyinput330,keyinput331,keyinput332,
keyinput333,keyinput334,keyinput335,keyinput336,keyinput337,keyinput338,keyinput339,keyinput340,keyinput341,keyinput342,
keyinput343,keyinput344,keyinput345,keyinput346,keyinput347,keyinput348,keyinput349,keyinput350,keyinput351,keyinput352,
keyinput353,keyinput354,keyinput355,keyinput356,keyinput357,keyinput358,keyinput359,keyinput360,keyinput361,keyinput362,
keyinput363,keyinput364,keyinput365,keyinput366,keyinput367,keyinput368,keyinput369,keyinput370,keyinput371,keyinput372,
keyinput373,keyinput374,keyinput375,keyinput376,keyinput377,keyinput378,keyinput379,keyinput380,keyinput381,keyinput382,
keyinput383,keyinput384,keyinput385,keyinput386,keyinput387);

input G1gat,G8gat,G13gat,G17gat,G26gat,G29gat,G36gat,G42gat,G51gat,
G55gat,G59gat,G68gat,G72gat,G73gat,G74gat,G75gat,G80gat,G85gat,G86gat,
G87gat,G88gat,G89gat,G90gat,G91gat,G96gat,G101gat,G106gat,G111gat,G116gat,
G121gat,G126gat,G130gat,G135gat,G138gat,G143gat,G146gat,G149gat,G152gat,G153gat,
G156gat,G159gat,G165gat,G171gat,G177gat,G183gat,G189gat,G195gat,G201gat,G207gat,
G210gat,G219gat,G228gat,G237gat,G246gat,G255gat,G259gat,G260gat,G261gat,G267gat,
G268gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,
keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,
keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,
keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,keyinput38,
keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,keyinput48,
keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,keyinput55,keyinput56,keyinput57,keyinput58,
keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,keyinput65,keyinput66,keyinput67,keyinput68,
keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,keyinput75,keyinput76,keyinput77,keyinput78,
keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,keyinput85,keyinput86,keyinput87,keyinput88,
keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,keyinput95,keyinput96,keyinput97,keyinput98,
keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,keyinput105,keyinput106,keyinput107,keyinput108,
keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,keyinput115,keyinput116,keyinput117,keyinput118,
keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,keyinput125,keyinput126,keyinput127,keyinput128,
keyinput129,keyinput130,keyinput131,keyinput132,keyinput133,keyinput134,keyinput135,keyinput136,keyinput137,keyinput138,
keyinput139,keyinput140,keyinput141,keyinput142,keyinput143,keyinput144,keyinput145,keyinput146,keyinput147,keyinput148,
keyinput149,keyinput150,keyinput151,keyinput152,keyinput153,keyinput154,keyinput155,keyinput156,keyinput157,keyinput158,
keyinput159,keyinput160,keyinput161,keyinput162,keyinput163,keyinput164,keyinput165,keyinput166,keyinput167,keyinput168,
keyinput169,keyinput170,keyinput171,keyinput172,keyinput173,keyinput174,keyinput175,keyinput176,keyinput177,keyinput178,
keyinput179,keyinput180,keyinput181,keyinput182,keyinput183,keyinput184,keyinput185,keyinput186,keyinput187,keyinput188,
keyinput189,keyinput190,keyinput191,keyinput192,keyinput193,keyinput194,keyinput195,keyinput196,keyinput197,keyinput198,
keyinput199,keyinput200,keyinput201,keyinput202,keyinput203,keyinput204,keyinput205,keyinput206,keyinput207,keyinput208,
keyinput209,keyinput210,keyinput211,keyinput212,keyinput213,keyinput214,keyinput215,keyinput216,keyinput217,keyinput218,
keyinput219,keyinput220,keyinput221,keyinput222,keyinput223,keyinput224,keyinput225,keyinput226,keyinput227,keyinput228,
keyinput229,keyinput230,keyinput231,keyinput232,keyinput233,keyinput234,keyinput235,keyinput236,keyinput237,keyinput238,
keyinput239,keyinput240,keyinput241,keyinput242,keyinput243,keyinput244,keyinput245,keyinput246,keyinput247,keyinput248,
keyinput249,keyinput250,keyinput251,keyinput252,keyinput253,keyinput254,keyinput255,keyinput256,keyinput257,keyinput258,
keyinput259,keyinput260,keyinput261,keyinput262,keyinput263,keyinput264,keyinput265,keyinput266,keyinput267,keyinput268,
keyinput269,keyinput270,keyinput271,keyinput272,keyinput273,keyinput274,keyinput275,keyinput276,keyinput277,keyinput278,
keyinput279,keyinput280,keyinput281,keyinput282,keyinput283,keyinput284,keyinput285,keyinput286,keyinput287,keyinput288,
keyinput289,keyinput290,keyinput291,keyinput292,keyinput293,keyinput294,keyinput295,keyinput296,keyinput297,keyinput298,
keyinput299,keyinput300,keyinput301,keyinput302,keyinput303,keyinput304,keyinput305,keyinput306,keyinput307,keyinput308,
keyinput309,keyinput310,keyinput311,keyinput312,keyinput313,keyinput314,keyinput315,keyinput316,keyinput317,keyinput318,
keyinput319,keyinput320,keyinput321,keyinput322,keyinput323,keyinput324,keyinput325,keyinput326,keyinput327,keyinput328,
keyinput329,keyinput330,keyinput331,keyinput332,keyinput333,keyinput334,keyinput335,keyinput336,keyinput337,keyinput338,
keyinput339,keyinput340,keyinput341,keyinput342,keyinput343,keyinput344,keyinput345,keyinput346,keyinput347,keyinput348,
keyinput349,keyinput350,keyinput351,keyinput352,keyinput353,keyinput354,keyinput355,keyinput356,keyinput357,keyinput358,
keyinput359,keyinput360,keyinput361,keyinput362,keyinput363,keyinput364,keyinput365,keyinput366,keyinput367,keyinput368,
keyinput369,keyinput370,keyinput371,keyinput372,keyinput373,keyinput374,keyinput375,keyinput376,keyinput377,keyinput378,
keyinput379,keyinput380,keyinput381,keyinput382,keyinput383,keyinput384,keyinput385,keyinput386,keyinput387;

output G388gat,G389gat,G390gat,G391gat,G418gat,G419gat,G420gat,G421gat,G422gat,
G423gat,G446gat,G447gat,G448gat,G449gat,G450gat,G767gat,G768gat,G850gat,G863gat,
G864gat,G865gat,G866gat,G874gat,G878gat,G879gat,G880gat;

wire G269gat,G270gat,G273gat,G276gat,G279gat,G280gat,G284gat,G285gat,G286gat,
G287gat,G290gat,G291gat,G292gat,G293gat,G294gat,G295gat,G296gat,G297gat,G298gat,
G301gat,G302gat,G303gat,G304gat,G305gat,G306gat,G307gat,G308gat,G309gat,G310gat,
G316gat,G317gat,G318gat,G319gat,G322gat,G323gat,G324gat,G325gat,G326gat,G327gat,
G328gat,G329gat,G330gat,G331gat,G332gat,G333gat,G334gat,G335gat,G336gat,G337gat,
G338gat,G339gat,G340gat,G341gat,G342gat,G343gat,G344gat,G345gat,G346gat,G347gat,
G348gat,G349gat,G350gat,G351gat,G352gat,G353gat,G354gat,G355gat,G356gat,G357gat,
G360gat,G363gat,G366gat,G369gat,G375gat,G376gat,G379gat,G382gat,G385gat,G392gat,
G393gat,G399gat,G400gat,G401gat,G402gat,G403gat,G404gat,G405gat,G406gat,G407gat,
G408gat,G409gat,G410gat,G411gat,G412gat,G413gat,G414gat,G415gat,G416gat,G417gat,
G424gat,G425gat,G426gat,G427gat,G432gat,G437gat,G442gat,G443gat,G444gat,G445gat,
G451gat,G460gat,G463gat,G466gat,G475gat,G476gat,G477gat,G478gat,G479gat,G480gat,
G481gat,G482gat,G483gat,G488gat,G489gat,G490gat,G491gat,G492gat,G495gat,G498gat,
G499gat,G500gat,G501gat,G502gat,G503gat,G504gat,G505gat,G506gat,G507gat,G508gat,
G509gat,G510gat,G511gat,G512gat,G513gat,G514gat,G515gat,G516gat,G517gat,G518gat,
G519gat,G520gat,G521gat,G522gat,G523gat,G524gat,G525gat,G526gat,G527gat,G528gat,
G529gat,G530gat,G533gat,G536gat,G537gat,G538gat,G539gat,G540gat,G541gat,G542gat,
G543gat,G544gat,G547gat,G550gat,G551gat,G552gat,G553gat,G557gat,G561gat,G565gat,
G569gat,G573gat,G577gat,G581gat,G585gat,G586gat,G587gat,G588gat,G589gat,G590gat,
G593gat,G596gat,G597gat,G600gat,G605gat,G606gat,G609gat,G615gat,G616gat,G619gat,
G624gat,G625gat,G628gat,G631gat,G632gat,G635gat,G640gat,G641gat,G644gat,G650gat,
G651gat,G654gat,G659gat,G660gat,G661gat,G662gat,G665gat,G669gat,G670gat,G673gat,
G677gat,G678gat,G682gat,G686gat,G687gat,G692gat,G696gat,G697gat,G700gat,G704gat,
G705gat,G708gat,G712gat,G713gat,G717gat,G721gat,G722gat,G727gat,G731gat,G732gat,
G733gat,G734gat,G735gat,G736gat,G737gat,G738gat,G739gat,G740gat,G741gat,G742gat,
G743gat,G744gat,G745gat,G746gat,G747gat,G748gat,G749gat,G750gat,G751gat,G752gat,
G753gat,G754gat,G755gat,G756gat,G757gat,G758gat,G759gat,G760gat,G761gat,G762gat,
G763gat,G764gat,G765gat,G766gat,G769gat,G770gat,G771gat,G772gat,G773gat,G777gat,
G778gat,G781gat,G782gat,G785gat,G786gat,G787gat,G788gat,G789gat,G790gat,G791gat,
G792gat,G793gat,G794gat,G795gat,G796gat,G802gat,G803gat,G804gat,G805gat,G806gat,
G807gat,G808gat,G809gat,G810gat,G811gat,G812gat,G813gat,G814gat,G815gat,G819gat,
G822gat,G825gat,G826gat,G827gat,G828gat,G829gat,G830gat,G831gat,G832gat,G833gat,
G834gat,G835gat,G836gat,G837gat,G838gat,G839gat,G840gat,G841gat,G842gat,G843gat,
G844gat,G845gat,G846gat,G847gat,G848gat,G849gat,G851gat,G852gat,G853gat,G854gat,
G855gat,G856gat,G857gat,G858gat,G859gat,G860gat,G861gat,G862gat,G867gat,G868gat,
G869gat,G870gat,G871gat,G872gat,G873gat,G875gat,G876gat,G877gat,muxed0,muxed1,
muxed2,muxed3,muxed4,muxed5,muxed6,muxed7,muxed8,muxed9,muxed10,muxed11,
muxed12,muxed13,muxed14,muxed15,muxed16,muxed17,muxed18,muxed19,muxed20,muxed21,
muxed22,muxed23,muxed24,muxed25,muxed26,muxed27,muxed28,muxed29,muxed30,muxed31,
muxed32,muxed33,muxed34,muxed35,muxed36,muxed37,muxed38,muxed39,muxed40,muxed41,
muxed42,muxed43,muxed44,muxed45,muxed46,muxed47,muxed48,muxed49,muxed50,muxed51,
muxed52,muxed53,muxed54,muxed55,muxed56,muxed57,muxed58,muxed59,muxed60,muxed61,
muxed62,muxed63,muxed64,muxed65,muxed66,muxed67,muxed68,muxed69,muxed70,muxed71,
muxed72,muxed73,muxed74,muxed75,muxed76,muxed77,muxed78,muxed79,muxed80,muxed81,
muxed82,muxed83,muxed84,muxed85,muxed86,muxed87,muxed88,muxed89,muxed90,muxed91,
muxed92,muxed93,muxed94,muxed95,muxed96,muxed97,muxed98,muxed99,muxed100,muxed101,
muxed102,muxed103,muxed104,muxed105,muxed106,muxed107,muxed108,muxed109,muxed110,muxed111,
muxed112,muxed113,muxed114,muxed115,muxed116,muxed117,muxed118,muxed119,muxed120,muxed121,
muxed122,muxed123,muxed124,muxed125,muxed126,muxed127,muxed128,muxed129,muxed130,muxed131,
muxed132,muxed133,muxed134,muxed135,muxed136,muxed137,muxed138,muxed139,muxed140,muxed141,
muxed142,muxed143,muxed144,muxed145,muxed146,muxed147,muxed148,muxed149,muxed150,muxed151,
muxed152,muxed153,muxed154,muxed155,muxed156,muxed157,muxed158,muxed159,muxed160,muxed161,
muxed162,muxed163,muxed164,muxed165,muxed166,muxed167,muxed168,muxed169,muxed170,muxed171,
muxed172,muxed173,muxed174,muxed175,muxed176,muxed177,muxed178,muxed179,muxed180,muxed181,
muxed182,muxed183,muxed184,muxed185,muxed186,muxed187,muxed188,muxed189,muxed190,muxed191,
muxed192,muxed193,muxed194,muxed195,muxed196,muxed197,muxed198,muxed199,muxed200,muxed201,
muxed202,muxed203,muxed204,muxed205,muxed206,muxed207,muxed208,muxed209,muxed210,muxed211,
muxed212,muxed213,muxed214,muxed215,muxed216,muxed217,muxed218,muxed219,muxed220,muxed221,
muxed222,muxed223,muxed224,muxed225,muxed226,muxed227,muxed228,muxed229,muxed230,muxed231,
muxed232,muxed233,muxed234,muxed235,muxed236,muxed237,muxed238,muxed239,muxed240,muxed241,
muxed242,muxed243,muxed244,muxed245,muxed246,muxed247,muxed248,muxed249,muxed250,muxed251,
muxed252,muxed253,muxed254,muxed255,muxed256,muxed257,muxed258,muxed259,muxed260,muxed261,
muxed262,muxed263,muxed264,muxed265,muxed266,muxed267,muxed268,muxed269,muxed270,muxed271,
muxed272,muxed273,muxed274,muxed275,muxed276,muxed277,muxed278,muxed279,muxed280,muxed281,
muxed282,muxed283,muxed284,muxed285,muxed286,muxed287,muxed288,muxed289,muxed290,muxed291,
muxed292,muxed293,muxed294,muxed295,muxed296,muxed297,muxed298,muxed299,muxed300,muxed301,
muxed302,muxed303,muxed304,muxed305,muxed306,muxed307,muxed308,muxed309,muxed310,muxed311,
muxed312,muxed313,muxed314,muxed315,muxed316,muxed317,muxed318,muxed319,muxed320,muxed321,
muxed322,muxed323,muxed324,muxed325,muxed326,muxed327,muxed328,muxed329,muxed330,muxed331,
muxed332,muxed333,muxed334,muxed335,muxed336,muxed337,muxed338,muxed339,muxed340,muxed341,
muxed342,muxed343,muxed344,muxed345,muxed346,muxed347,muxed348,muxed349,muxed350,muxed351,
muxed352,muxed353,muxed354,muxed355,muxed356,muxed357,muxed358,muxed359,muxed360,muxed361,
muxed362,muxed363,muxed364,muxed365,muxed366,muxed367,muxed368,muxed369,muxed370,muxed371,
muxed372,muxed373,muxed374,muxed375,muxed376,muxed377,muxed378,muxed379,muxed380,muxed381,
muxed382,muxed383,muxed384,muxed385,muxed386,muxed387;
nand gate_0(G269gat,G1gat,G8gat,G13gat,G17gat);
nand gate_1(G270gat,G1gat,G26gat,G13gat,G17gat);
and gate_2(G273gat,G29gat,G36gat,G42gat);
and gate_3(G276gat,G1gat,G26gat,muxed270);
nand gate_4(G279gat,G1gat,G8gat,muxed270,G17gat);
nand gate_5(G280gat,G1gat,G8gat,G13gat,G55gat);
nand gate_6(G284gat,G59gat,G42gat,G68gat,G72gat);
nand gate_7(G285gat,G29gat,G68gat);
nand gate_8(G286gat,G59gat,G68gat,G74gat);
and gate_9(G287gat,G29gat,G75gat,G80gat);
and gate_10(G290gat,G29gat,G75gat,G42gat);
and gate_11(G291gat,G29gat,G36gat,G80gat);
and gate_12(G292gat,G29gat,G36gat,G42gat);
and gate_13(G293gat,G59gat,G75gat,G80gat);
and gate_14(G294gat,G59gat,G75gat,G42gat);
and gate_15(G295gat,G59gat,G36gat,G80gat);
and gate_16(G296gat,G59gat,G36gat,G42gat);
and gate_17(G297gat,G85gat,G86gat);
or gate_18(G298gat,G87gat,G88gat);
nand gate_19(G301gat,G91gat,G96gat);
or gate_20(G302gat,G91gat,G96gat);
nand gate_21(G303gat,G101gat,G106gat);
or gate_22(G304gat,G101gat,G106gat);
nand gate_23(G305gat,G111gat,G116gat);
or gate_24(G306gat,G111gat,G116gat);
nand gate_25(G307gat,muxed52,G126gat);
or gate_26(G308gat,muxed52,G126gat);
and gate_27(G309gat,G8gat,G138gat);
not gate_28(G310gat,G268gat);
and gate_29(G316gat,muxed270,G138gat);
and gate_30(G317gat,G17gat,G138gat);
and gate_31(G318gat,G152gat,G138gat);
nand gate_32(G319gat,G59gat,G156gat);
nor gate_33(G322gat,G17gat,G42gat);
and gate_34(G323gat,G17gat,G42gat);
nand gate_35(G324gat,G159gat,G165gat);
or gate_36(G325gat,G159gat,G165gat);
nand gate_37(G326gat,G171gat,G177gat);
or gate_38(G327gat,G171gat,G177gat);
nand gate_39(G328gat,G183gat,G189gat);
or gate_40(G329gat,G183gat,G189gat);
nand gate_41(G330gat,G195gat,G201gat);
or gate_42(G331gat,G195gat,G201gat);
and gate_43(G332gat,G210gat,G91gat);
and gate_44(G333gat,G210gat,G96gat);
and gate_45(G334gat,G210gat,G101gat);
and gate_46(G335gat,G210gat,G106gat);
and gate_47(G336gat,G210gat,G111gat);
and gate_48(G337gat,G255gat,G259gat);
and gate_49(G338gat,G210gat,G116gat);
and gate_50(G339gat,G255gat,G260gat);
and gate_51(G340gat,G210gat,muxed52);
and gate_52(G341gat,G255gat,G267gat);
not gate_53(G342gat,G269gat);
not gate_54(G343gat,G273gat);
or gate_55(G344gat,G270gat,G273gat);
not gate_56(G345gat,muxed76);
not gate_57(G346gat,muxed76);
not gate_58(G347gat,G279gat);
nor gate_59(G348gat,G280gat,G284gat);
or gate_60(G349gat,G280gat,G285gat);
or gate_61(G350gat,G280gat,G286gat);
not gate_62(G351gat,muxed246);
not gate_63(G352gat,G294gat);
not gate_64(G353gat,muxed352);
not gate_65(G354gat,G296gat);
nand gate_66(G355gat,G89gat,muxed237);
and gate_67(G356gat,G90gat,muxed237);
nand gate_68(G357gat,muxed111,G302gat);
nand gate_69(G360gat,muxed320,G304gat);
nand gate_70(G363gat,G305gat,G306gat);
nand gate_71(G366gat,G307gat,G308gat);
not gate_72(G369gat,G310gat);
nor gate_73(G375gat,G322gat,G323gat);
nand gate_74(G376gat,muxed188,G325gat);
nand gate_75(G379gat,G326gat,G327gat);
nand gate_76(G382gat,G328gat,G329gat);
nand gate_77(G385gat,G330gat,G331gat);
buf gate_78(G388gat,G290gat);
buf gate_79(G389gat,G291gat);
buf gate_80(G390gat,G292gat);
buf gate_81(G391gat,G297gat);
or gate_82(G392gat,G270gat,G343gat);
not gate_83(G393gat,muxed97);
not gate_84(G399gat,G346gat);
and gate_85(G400gat,G348gat,G73gat);
not gate_86(G401gat,muxed51);
not gate_87(G402gat,G350gat);
not gate_88(G403gat,G355gat);
not gate_89(G404gat,G357gat);
not gate_90(G405gat,muxed319);
and gate_91(G406gat,G357gat,muxed319);
not gate_92(G407gat,muxed196);
not gate_93(G408gat,G366gat);
and gate_94(G409gat,muxed196,G366gat);
nand gate_95(G410gat,G347gat,G352gat);
not gate_96(G411gat,muxed156);
not gate_97(G412gat,G379gat);
and gate_98(G413gat,muxed156,G379gat);
not gate_99(G414gat,G382gat);
not gate_100(G415gat,muxed94);
and gate_101(G416gat,G382gat,muxed94);
and gate_102(G417gat,G210gat,muxed338);
buf gate_103(G418gat,G342gat);
buf gate_104(G419gat,G344gat);
buf gate_105(G420gat,G351gat);
buf gate_106(G421gat,muxed174);
buf gate_107(G422gat,G354gat);
buf gate_108(G423gat,G356gat);
not gate_109(G424gat,muxed151);
and gate_110(G425gat,muxed9,G405gat);
and gate_111(G426gat,G407gat,G408gat);
and gate_112(G427gat,G319gat,muxed315,G55gat);
and gate_113(G432gat,muxed315,G17gat,G287gat);
nand gate_114(G437gat,muxed315,G287gat,G55gat);
nand gate_115(G442gat,G375gat,G59gat,G156gat,muxed315);
nand gate_116(G443gat,muxed315,G319gat,G17gat);
and gate_117(G444gat,G411gat,G412gat);
and gate_118(G445gat,G414gat,muxed265);
buf gate_119(G446gat,G392gat);
buf gate_120(G447gat,G399gat);
buf gate_121(G448gat,G401gat);
buf gate_122(G449gat,G402gat);
buf gate_123(G450gat,G403gat);
not gate_124(G451gat,G424gat);
nor gate_125(G460gat,muxed317,G425gat);
nor gate_126(G463gat,G409gat,G426gat);
nand gate_127(G466gat,G442gat,muxed155);
and gate_128(G475gat,G143gat,G427gat);
and gate_129(G476gat,G310gat,muxed354);
and gate_130(G477gat,G146gat,G427gat);
and gate_131(G478gat,G310gat,muxed354);
and gate_132(G479gat,G149gat,G427gat);
and gate_133(G480gat,G310gat,muxed354);
and gate_134(G481gat,G153gat,G427gat);
and gate_135(G482gat,G310gat,muxed354);
nand gate_136(G483gat,muxed193,G1gat);
or gate_137(G488gat,muxed338,muxed337);
or gate_138(G489gat,muxed338,muxed337);
or gate_139(G490gat,muxed338,muxed337);
or gate_140(G491gat,muxed338,muxed337);
nor gate_141(G492gat,muxed153,G444gat);
nor gate_142(G495gat,muxed59,G445gat);
nand gate_143(G498gat,G130gat,muxed22);
or gate_144(G499gat,G130gat,muxed22);
nand gate_145(G500gat,G463gat,G135gat);
or gate_146(G501gat,G463gat,G135gat);
and gate_147(G502gat,G91gat,muxed165);
nor gate_148(G503gat,G475gat,G476gat);
and gate_149(G504gat,G96gat,muxed165);
nor gate_150(G505gat,G477gat,muxed136);
and gate_151(G506gat,G101gat,muxed165);
nor gate_152(G507gat,G479gat,G480gat);
and gate_153(G508gat,G106gat,muxed165);
nor gate_154(G509gat,muxed259,G482gat);
and gate_155(G510gat,G143gat,G483gat);
and gate_156(G511gat,G111gat,muxed165);
and gate_157(G512gat,G146gat,G483gat);
and gate_158(G513gat,G116gat,muxed165);
and gate_159(G514gat,G149gat,G483gat);
and gate_160(G515gat,muxed52,muxed165);
and gate_161(G516gat,G153gat,G483gat);
and gate_162(G517gat,G126gat,muxed165);
nand gate_163(G518gat,G130gat,G492gat);
or gate_164(G519gat,G130gat,G492gat);
nand gate_165(G520gat,muxed37,G207gat);
or gate_166(G521gat,muxed37,G207gat);
and gate_167(G522gat,G451gat,G159gat);
and gate_168(G523gat,G451gat,G165gat);
and gate_169(G524gat,G451gat,G171gat);
and gate_170(G525gat,G451gat,G177gat);
and gate_171(G526gat,G451gat,G183gat);
nand gate_172(G527gat,G451gat,G189gat);
nand gate_173(G528gat,G451gat,G195gat);
nand gate_174(G529gat,G451gat,G201gat);
nand gate_175(G530gat,muxed261,G499gat);
nand gate_176(G533gat,muxed332,G501gat);
nor gate_177(G536gat,G309gat,G502gat);
nor gate_178(G537gat,muxed293,G504gat);
nor gate_179(G538gat,muxed167,G506gat);
nor gate_180(G539gat,G318gat,G508gat);
nor gate_181(G540gat,G510gat,muxed206);
nor gate_182(G541gat,G512gat,G513gat);
nor gate_183(G542gat,G514gat,muxed335);
nor gate_184(G543gat,G516gat,G517gat);
nand gate_185(G544gat,G518gat,G519gat);
nand gate_186(G547gat,muxed140,muxed35);
not gate_187(G550gat,muxed260);
not gate_188(G551gat,muxed369);
and gate_189(G552gat,muxed260,muxed369);
nand gate_190(G553gat,G536gat,G503gat);
nand gate_191(G557gat,muxed159,G505gat);
nand gate_192(G561gat,G538gat,muxed255);
nand gate_193(G565gat,G539gat,G509gat);
nand gate_194(G569gat,muxed360,muxed229);
nand gate_195(G573gat,muxed84,G541gat);
nand gate_196(G577gat,muxed192,muxed72);
nand gate_197(G581gat,muxed248,G543gat);
not gate_198(G585gat,G544gat);
not gate_199(G586gat,muxed321);
and gate_200(G587gat,G544gat,muxed321);
and gate_201(G588gat,G550gat,G551gat);
and gate_202(G589gat,muxed182,G586gat);
nand gate_203(G590gat,G553gat,G159gat);
or gate_204(G593gat,G553gat,G159gat);
and gate_205(G596gat,G246gat,G553gat);
nand gate_206(G597gat,muxed158,G165gat);
or gate_207(G600gat,muxed158,G165gat);
and gate_208(G605gat,G246gat,muxed158);
nand gate_209(G606gat,G561gat,G171gat);
or gate_210(G609gat,G561gat,G171gat);
and gate_211(G615gat,G246gat,G561gat);
nand gate_212(G616gat,muxed238,G177gat);
or gate_213(G619gat,muxed238,G177gat);
and gate_214(G624gat,G246gat,muxed238);
nand gate_215(G625gat,muxed256,G183gat);
or gate_216(G628gat,muxed256,G183gat);
and gate_217(G631gat,G246gat,muxed256);
nand gate_218(G632gat,muxed24,G189gat);
or gate_219(G635gat,muxed24,G189gat);
and gate_220(G640gat,G246gat,muxed24);
nand gate_221(G641gat,muxed127,G195gat);
or gate_222(G644gat,muxed127,G195gat);
and gate_223(G650gat,G246gat,muxed127);
nand gate_224(G651gat,G581gat,G201gat);
or gate_225(G654gat,G581gat,G201gat);
and gate_226(G659gat,G246gat,G581gat);
nor gate_227(G660gat,muxed258,G588gat);
nor gate_228(G661gat,muxed32,muxed181);
not gate_229(G662gat,G590gat);
and gate_230(G665gat,muxed163,G590gat);
nor gate_231(G669gat,muxed93,G522gat);
not gate_232(G670gat,G597gat);
and gate_233(G673gat,muxed297,G597gat);
nor gate_234(G677gat,muxed157,G523gat);
not gate_235(G678gat,G606gat);
and gate_236(G682gat,G609gat,G606gat);
nor gate_237(G686gat,G615gat,G524gat);
not gate_238(G687gat,G616gat);
and gate_239(G692gat,G619gat,G616gat);
nor gate_240(G696gat,muxed233,G525gat);
not gate_241(G697gat,muxed230);
and gate_242(G700gat,G628gat,muxed230);
nor gate_243(G704gat,muxed201,G526gat);
not gate_244(G705gat,G632gat);
and gate_245(G708gat,muxed23,G632gat);
nor gate_246(G712gat,G337gat,G640gat);
not gate_247(G713gat,muxed200);
and gate_248(G717gat,G644gat,muxed200);
nor gate_249(G721gat,muxed305,G650gat);
not gate_250(G722gat,G651gat);
and gate_251(G727gat,muxed232,G651gat);
nor gate_252(G731gat,G341gat,G659gat);
nand gate_253(G732gat,muxed232,G261gat);
nand gate_254(G733gat,G644gat,muxed232,G261gat);
nand gate_255(G734gat,muxed23,G644gat,muxed232,G261gat);
not gate_256(G735gat,G662gat);
and gate_257(G736gat,G228gat,muxed162);
and gate_258(G737gat,muxed27,G662gat);
not gate_259(G738gat,muxed362);
and gate_260(G739gat,G228gat,G673gat);
and gate_261(G740gat,muxed27,muxed362);
not gate_262(G741gat,muxed114);
and gate_263(G742gat,G228gat,G682gat);
and gate_264(G743gat,muxed27,muxed114);
not gate_265(G744gat,muxed33);
and gate_266(G745gat,G228gat,G692gat);
and gate_267(G746gat,muxed27,muxed33);
not gate_268(G747gat,G697gat);
and gate_269(G748gat,G228gat,G700gat);
and gate_270(G749gat,muxed27,G697gat);
not gate_271(G750gat,G705gat);
and gate_272(G751gat,G228gat,muxed26);
and gate_273(G752gat,muxed27,G705gat);
not gate_274(G753gat,G713gat);
and gate_275(G754gat,G228gat,G717gat);
and gate_276(G755gat,muxed27,G713gat);
not gate_277(G756gat,muxed205);
nor gate_278(G757gat,G727gat,G261gat);
and gate_279(G758gat,G727gat,G261gat);
and gate_280(G759gat,G228gat,G727gat);
and gate_281(G760gat,muxed27,muxed205);
nand gate_282(G761gat,G644gat,muxed205);
nand gate_283(G762gat,muxed23,G713gat);
nand gate_284(G763gat,muxed23,G644gat,muxed205);
nand gate_285(G764gat,G609gat,muxed33);
nand gate_286(G765gat,muxed297,muxed114);
nand gate_287(G766gat,muxed297,G609gat,muxed33);
buf gate_288(G767gat,muxed257);
buf gate_289(G768gat,muxed30);
nor gate_290(G769gat,G736gat,G737gat);
nor gate_291(G770gat,G739gat,G740gat);
nor gate_292(G771gat,G742gat,G743gat);
nor gate_293(G772gat,G745gat,G746gat);
nand gate_294(G773gat,muxed173,G762gat,muxed21,muxed231);
nor gate_295(G777gat,G748gat,G749gat);
nand gate_296(G778gat,G753gat,muxed175,G733gat);
nor gate_297(G781gat,muxed247,muxed50);
nand gate_298(G782gat,muxed180,muxed148);
nor gate_299(G785gat,muxed197,G755gat);
nor gate_300(G786gat,G757gat,G758gat);
nor gate_301(G787gat,muxed235,G760gat);
nor gate_302(G788gat,G700gat,muxed20);
and gate_303(G789gat,G700gat,muxed20);
nor gate_304(G790gat,muxed26,G778gat);
and gate_305(G791gat,muxed26,G778gat);
nor gate_306(G792gat,G717gat,muxed366);
and gate_307(G793gat,G717gat,muxed366);
and gate_308(G794gat,G219gat,G786gat);
nand gate_309(G795gat,G628gat,muxed20);
nand gate_310(G796gat,muxed85,G747gat);
nor gate_311(G802gat,muxed281,G789gat);
nor gate_312(G803gat,G790gat,G791gat);
nor gate_313(G804gat,G792gat,muxed209);
nor gate_314(G805gat,muxed36,G794gat);
nor gate_315(G806gat,G692gat,muxed80);
and gate_316(G807gat,G692gat,muxed80);
and gate_317(G808gat,G219gat,muxed279);
and gate_318(G809gat,G219gat,G803gat);
and gate_319(G810gat,G219gat,muxed141);
nand gate_320(G811gat,G805gat,G787gat,G731gat,muxed149);
nand gate_321(G812gat,G619gat,muxed80);
nand gate_322(G813gat,G609gat,G619gat,muxed80);
nand gate_323(G814gat,muxed297,G609gat,G619gat,muxed80);
nand gate_324(G815gat,muxed385,G765gat,muxed56,muxed118);
nand gate_325(G819gat,G741gat,G764gat,G813gat);
nand gate_326(G822gat,G744gat,G812gat);
nor gate_327(G825gat,G806gat,G807gat);
nor gate_328(G826gat,G335gat,muxed277);
nor gate_329(G827gat,muxed98,G809gat);
nor gate_330(G828gat,G338gat,muxed137);
not gate_331(G829gat,muxed189);
nor gate_332(G830gat,muxed162,muxed68);
and gate_333(G831gat,muxed162,muxed68);
nor gate_334(G832gat,G673gat,G819gat);
and gate_335(G833gat,G673gat,G819gat);
nor gate_336(G834gat,G682gat,G822gat);
and gate_337(G835gat,G682gat,G822gat);
and gate_338(G836gat,G219gat,G825gat);
nand gate_339(G837gat,muxed171,G777gat,muxed199);
nand gate_340(G838gat,muxed75,muxed267,G712gat,G527gat);
nand gate_341(G839gat,muxed135,muxed342,muxed19,G528gat);
not gate_342(G840gat,G829gat);
nand gate_343(G841gat,muxed68,muxed163);
nor gate_344(G842gat,muxed264,muxed12);
nor gate_345(G843gat,G832gat,G833gat);
nor gate_346(G844gat,G834gat,G835gat);
nor gate_347(G845gat,G334gat,G836gat);
not gate_348(G846gat,muxed195);
not gate_349(G847gat,muxed324);
not gate_350(G848gat,muxed218);
and gate_351(G849gat,G735gat,G841gat);
buf gate_352(G850gat,G840gat);
and gate_353(G851gat,G219gat,muxed371);
and gate_354(G852gat,G219gat,G843gat);
and gate_355(G853gat,G219gat,G844gat);
nand gate_356(G854gat,G845gat,G772gat,G696gat);
not gate_357(G855gat,muxed194);
not gate_358(G856gat,muxed312);
not gate_359(G857gat,muxed240);
not gate_360(G858gat,G849gat);
nor gate_361(G859gat,G417gat,muxed177);
nor gate_362(G860gat,G332gat,G852gat);
nor gate_363(G861gat,G333gat,G853gat);
not gate_364(G862gat,G854gat);
buf gate_365(G863gat,G855gat);
buf gate_366(G864gat,muxed123);
buf gate_367(G865gat,G857gat);
buf gate_368(G866gat,G858gat);
nand gate_369(G867gat,muxed53,G769gat,G669gat);
nand gate_370(G868gat,G860gat,G770gat,muxed39);
nand gate_371(G869gat,G861gat,G771gat,G686gat);
not gate_372(G870gat,G862gat);
not gate_373(G871gat,muxed4);
not gate_374(G872gat,G868gat);
not gate_375(G873gat,muxed311);
buf gate_376(G874gat,G870gat);
not gate_377(G875gat,muxed2);
not gate_378(G876gat,G872gat);
not gate_379(G877gat,G873gat);
buf gate_380(G878gat,muxed1);
buf gate_381(G879gat,G876gat);
buf gate_382(G880gat,G877gat);
assign muxed0 = keyinput0 ? G369gat : muxed1;
assign muxed1 = keyinput1 ? muxed278 : G544gat;
assign muxed2 = keyinput2 ? G871gat : G845gat;
assign muxed3 = keyinput3 ? muxed283 : G871gat;
assign muxed4 = keyinput4 ? muxed207 : muxed293;
assign muxed5 = keyinput5 ? muxed146 : muxed207;
assign muxed6 = keyinput6 ? muxed176 : muxed369;
assign muxed7 = keyinput7 ? G353gat : muxed176;
assign muxed8 = keyinput8 ? G851gat : muxed181;
assign muxed9 = keyinput9 ? G404gat : G851gat;
assign muxed10 = keyinput10 ? muxed263 : muxed20;
assign muxed11 = keyinput11 ? muxed117 : muxed263;
assign muxed12 = keyinput12 ? muxed65 : G409gat;
assign muxed13 = keyinput13 ? muxed106 : muxed65;
assign muxed14 = keyinput14 ? muxed43 : muxed127;
assign muxed15 = keyinput15 ? muxed78 : muxed153;
assign muxed16 = keyinput16 ? G766gat : muxed78;
assign muxed17 = keyinput17 ? muxed83 : muxed267;
assign muxed18 = keyinput18 ? G795gat : muxed165;
assign muxed19 = keyinput19 ? G721gat : G795gat;
assign muxed20 = keyinput20 ? G773gat : G343gat;
assign muxed21 = keyinput21 ? muxed183 : G334gat;
assign muxed22 = keyinput22 ? muxed316 : muxed183;
assign muxed23 = keyinput23 ? G635gat : G757gat;
assign muxed24 = keyinput24 ? G573gat : G290gat;
assign muxed25 = keyinput25 ? muxed250 : G697gat;
assign muxed26 = keyinput26 ? G708gat : muxed250;
assign muxed27 = keyinput27 ? G237gat : muxed28;
assign muxed28 = keyinput28 ? G768gat : muxed167;
assign muxed29 = keyinput29 ? muxed122 : G768gat;
assign muxed30 = keyinput30 ? G661gat : G375gat;
assign muxed31 = keyinput31 ? muxed239 : G661gat;
assign muxed32 = keyinput32 ? G587gat : G286gat;
assign muxed33 = keyinput33 ? G687gat : G587gat;
assign muxed34 = keyinput34 ? G547gat : G426gat;
assign muxed35 = keyinput35 ? muxed107 : muxed26;
assign muxed36 = keyinput36 ? G340gat : muxed107;
assign muxed37 = keyinput37 ? muxed350 : muxed2;
assign muxed38 = keyinput38 ? muxed91 : muxed369;
assign muxed39 = keyinput39 ? G677gat : muxed91;
assign muxed40 = keyinput40 ? muxed103 : muxed362;
assign muxed41 = keyinput41 ? muxed66 : G851gat;
assign muxed42 = keyinput42 ? muxed69 : G748gat;
assign muxed43 = keyinput43 ? muxed115 : G794gat;
assign muxed44 = keyinput44 ? muxed64 : muxed115;
assign muxed45 = keyinput45 ? muxed77 : muxed350;
assign muxed46 = keyinput46 ? muxed185 : muxed77;
assign muxed47 = keyinput47 ? muxed336 : muxed371;
assign muxed48 = keyinput48 ? muxed81 : G644gat;
assign muxed49 = keyinput49 ? muxed374 : G753gat;
assign muxed50 = keyinput50 ? muxed214 : G765gat;
assign muxed51 = keyinput51 ? G349gat : muxed214;
assign muxed52 = keyinput52 ? G121gat : muxed53;
assign muxed53 = keyinput53 ? muxed6 : muxed265;
assign muxed54 = keyinput54 ? muxed113 : muxed305;
assign muxed55 = keyinput55 ? muxed116 : G354gat;
assign muxed56 = keyinput56 ? muxed212 : G547gat;
assign muxed57 = keyinput57 ? muxed341 : muxed212;
assign muxed58 = keyinput58 ? G495gat : muxed218;
assign muxed59 = keyinput59 ? muxed109 : muxed336;
assign muxed60 = keyinput60 ? G410gat : muxed109;
assign muxed61 = keyinput61 ? muxed346 : G651gat;
assign muxed62 = keyinput62 ? muxed101 : muxed193;
assign muxed63 = keyinput63 ? muxed105 : G692gat;
assign muxed64 = keyinput64 ? muxed331 : muxed105;
assign muxed65 = keyinput65 ? muxed41 : G417gat;
assign muxed66 = keyinput66 ? muxed217 : muxed385;
assign muxed67 = keyinput67 ? muxed381 : muxed217;
assign muxed68 = keyinput68 ? muxed42 : G586gat;
assign muxed69 = keyinput69 ? muxed126 : G697gat;
assign muxed70 = keyinput70 ? muxed274 : muxed126;
assign muxed71 = keyinput71 ? muxed128 : G509gat;
assign muxed72 = keyinput72 ? muxed334 : G807gat;
assign muxed73 = keyinput73 ? G500gat : muxed334;
assign muxed74 = keyinput74 ? G515gat : muxed337;
assign muxed75 = keyinput75 ? G827gat : G515gat;
assign muxed76 = keyinput76 ? G276gat : muxed77;
assign muxed77 = keyinput77 ? muxed16 : G342gat;
assign muxed78 = keyinput78 ? muxed47 : G310gat;
assign muxed79 = keyinput79 ? muxed329 : G536gat;
assign muxed80 = keyinput80 ? muxed48 : G845gat;
assign muxed81 = keyinput81 ? muxed266 : G334gat;
assign muxed82 = keyinput82 ? G830gat : muxed266;
assign muxed83 = keyinput83 ? G796gat : G424gat;
assign muxed84 = keyinput84 ? muxed25 : G796gat;
assign muxed85 = keyinput85 ? muxed358 : G697gat;
assign muxed86 = keyinput86 ? G593gat : muxed358;
assign muxed87 = keyinput87 ? muxed166 : muxed123;
assign muxed88 = keyinput88 ? muxed108 : muxed312;
assign muxed89 = keyinput89 ? G385gat : muxed108;
assign muxed90 = keyinput90 ? muxed292 : G581gat;
assign muxed91 = keyinput91 ? muxed61 : G337gat;
assign muxed92 = keyinput92 ? G416gat : muxed329;
assign muxed93 = keyinput93 ? G596gat : G416gat;
assign muxed94 = keyinput94 ? muxed190 : muxed149;
assign muxed95 = keyinput95 ? G443gat : muxed194;
assign muxed96 = keyinput96 ? muxed102 : muxed140;
assign muxed97 = keyinput97 ? G345gat : G480gat;
assign muxed98 = keyinput98 ? G336gat : G345gat;
assign muxed99 = keyinput99 ? G324gat : muxed190;
assign muxed100 = keyinput100 ? muxed191 : muxed247;
assign muxed101 = keyinput101 ? muxed40 : G740gat;
assign muxed102 = keyinput102 ? G393gat : muxed40;
assign muxed103 = keyinput103 ? muxed63 : muxed305;
assign muxed104 = keyinput104 ? G600gat : muxed63;
assign muxed105 = keyinput105 ? muxed13 : muxed235;
assign muxed106 = keyinput106 ? muxed372 : muxed68;
assign muxed107 = keyinput107 ? G521gat : muxed372;
assign muxed108 = keyinput108 ? muxed60 : muxed115;
assign muxed109 = keyinput109 ? muxed90 : G477gat;
assign muxed110 = keyinput110 ? muxed38 : G843gat;
assign muxed111 = keyinput111 ? muxed344 : muxed38;
assign muxed112 = keyinput112 ? muxed54 : muxed372;
assign muxed113 = keyinput113 ? muxed44 : G765gat;
assign muxed114 = keyinput114 ? G678gat : muxed44;
assign muxed115 = keyinput115 ? muxed55 : G319gat;
assign muxed116 = keyinput116 ? G815gat : G309gat;
assign muxed117 = keyinput117 ? G498gat : G815gat;
assign muxed118 = keyinput118 ? muxed152 : muxed41;
assign muxed119 = keyinput119 ? G400gat : muxed152;
assign muxed120 = keyinput120 ? muxed154 : G509gat;
assign muxed121 = keyinput121 ? muxed29 : muxed157;
assign muxed122 = keyinput122 ? muxed287 : G335gat;
assign muxed123 = keyinput123 ? muxed387 : muxed287;
assign muxed124 = keyinput124 ? G654gat : muxed233;
assign muxed125 = keyinput125 ? muxed234 : G640gat;
assign muxed126 = keyinput126 ? muxed14 : G553gat;
assign muxed127 = keyinput127 ? muxed71 : muxed240;
assign muxed128 = keyinput128 ? G577gat : muxed90;
assign muxed129 = keyinput129 ? muxed386 : G577gat;
assign muxed130 = keyinput130 ? muxed275 : G402gat;
assign muxed131 = keyinput131 ? muxed143 : muxed275;
assign muxed132 = keyinput132 ? muxed213 : G870gat;
assign muxed133 = keyinput133 ? muxed353 : muxed362;
assign muxed134 = keyinput134 ? muxed219 : G279gat;
assign muxed135 = keyinput135 ? G828gat : muxed113;
assign muxed136 = keyinput136 ? G478gat : G828gat;
assign muxed137 = keyinput137 ? muxed184 : G586gat;
assign muxed138 = keyinput138 ? G585gat : muxed184;
assign muxed139 = keyinput139 ? G810gat : muxed287;
assign muxed140 = keyinput140 ? G520gat : G810gat;
assign muxed141 = keyinput141 ? muxed208 : muxed205;
assign muxed142 = keyinput142 ? G511gat : muxed208;
assign muxed143 = keyinput143 ? muxed363 : G778gat;
assign muxed144 = keyinput144 ? muxed104 : muxed363;
assign muxed145 = keyinput145 ? muxed222 : muxed369;
assign muxed146 = keyinput146 ? G782gat : G845gat;
assign muxed147 = keyinput147 ? G722gat : G782gat;
assign muxed148 = keyinput148 ? muxed377 : muxed26;
assign muxed149 = keyinput149 ? G529gat : muxed377;
assign muxed150 = keyinput150 ? G838gat : muxed151;
assign muxed151 = keyinput151 ? muxed348 : muxed51;
assign muxed152 = keyinput152 ? muxed15 : G790gat;
assign muxed153 = keyinput153 ? muxed120 : G762gat;
assign muxed154 = keyinput154 ? G413gat : muxed344;
assign muxed155 = keyinput155 ? muxed168 : G413gat;
assign muxed156 = keyinput156 ? muxed121 : muxed65;
assign muxed157 = keyinput157 ? G605gat : muxed115;
assign muxed158 = keyinput158 ? G557gat : G606gat;
assign muxed159 = keyinput159 ? muxed378 : muxed52;
assign muxed160 = keyinput160 ? muxed179 : muxed378;
assign muxed161 = keyinput161 ? G831gat : muxed246;
assign muxed162 = keyinput162 ? G665gat : muxed127;
assign muxed163 = keyinput163 ? muxed355 : G877gat;
assign muxed164 = keyinput164 ? muxed18 : G351gat;
assign muxed165 = keyinput165 ? muxed87 : muxed98;
assign muxed166 = keyinput166 ? G466gat : G748gat;
assign muxed167 = keyinput167 ? G317gat : G466gat;
assign muxed168 = keyinput168 ? muxed307 : G677gat;
assign muxed169 = keyinput169 ? G788gat : muxed307;
assign muxed170 = keyinput170 ? muxed313 : G851gat;
assign muxed171 = keyinput171 ? muxed276 : muxed172;
assign muxed172 = keyinput172 ? G421gat : G868gat;
assign muxed173 = keyinput173 ? G750gat : G421gat;
assign muxed174 = keyinput174 ? muxed7 : muxed168;
assign muxed175 = keyinput175 ? G761gat : muxed7;
assign muxed176 = keyinput176 ? G859gat : G834gat;
assign muxed177 = keyinput177 ? muxed375 : muxed84;
assign muxed178 = keyinput178 ? muxed244 : muxed375;
assign muxed179 = keyinput179 ? muxed8 : G713gat;
assign muxed180 = keyinput180 ? G756gat : muxed8;
assign muxed181 = keyinput181 ? G589gat : G515gat;
assign muxed182 = keyinput182 ? muxed138 : muxed108;
assign muxed183 = keyinput183 ? G763gat : muxed138;
assign muxed184 = keyinput184 ? muxed46 : G763gat;
assign muxed185 = keyinput185 ? muxed286 : G692gat;
assign muxed186 = keyinput186 ? muxed310 : muxed286;
assign muxed187 = keyinput187 ? muxed288 : muxed46;
assign muxed188 = keyinput188 ? muxed99 : G369gat;
assign muxed189 = keyinput189 ? G811gat : muxed99;
assign muxed190 = keyinput190 ? muxed357 : G399gat;
assign muxed191 = keyinput191 ? muxed309 : G737gat;
assign muxed192 = keyinput192 ? muxed130 : muxed309;
assign muxed193 = keyinput193 ? muxed95 : muxed25;
assign muxed194 = keyinput194 ? G846gat : G758gat;
assign muxed195 = keyinput195 ? muxed198 : G355gat;
assign muxed196 = keyinput196 ? G363gat : muxed198;
assign muxed197 = keyinput197 ? G754gat : muxed198;
assign muxed198 = keyinput198 ? G837gat : G306gat;
assign muxed199 = keyinput199 ? G704gat : muxed235;
assign muxed200 = keyinput200 ? G641gat : G704gat;
assign muxed201 = keyinput201 ? muxed280 : G756gat;
assign muxed202 = keyinput202 ? G489gat : muxed280;
assign muxed203 = keyinput203 ? muxed227 : G597gat;
assign muxed204 = keyinput204 ? G540gat : muxed231;
assign muxed205 = keyinput205 ? muxed147 : G540gat;
assign muxed206 = keyinput206 ? muxed142 : G327gat;
assign muxed207 = keyinput207 ? G867gat : muxed142;
assign muxed208 = keyinput208 ? G804gat : muxed111;
assign muxed209 = keyinput209 ? muxed272 : muxed138;
assign muxed210 = keyinput210 ? G565gat : muxed272;
assign muxed211 = keyinput211 ? muxed243 : G516gat;
assign muxed212 = keyinput212 ? muxed132 : muxed76;
assign muxed213 = keyinput213 ? muxed349 : G749gat;
assign muxed214 = keyinput214 ? G752gat : muxed349;
assign muxed215 = keyinput215 ? muxed351 : G756gat;
assign muxed216 = keyinput216 ? muxed58 : muxed355;
assign muxed217 = keyinput217 ? muxed161 : muxed58;
assign muxed218 = keyinput218 ? muxed368 : G565gat;
assign muxed219 = keyinput219 ? muxed339 : G290gat;
assign muxed220 = keyinput220 ? muxed356 : muxed339;
assign muxed221 = keyinput221 ? G785gat : muxed344;
assign muxed222 = keyinput222 ? muxed5 : G785gat;
assign muxed223 = keyinput223 ? muxed0 : muxed250;
assign muxed224 = keyinput224 ? muxed251 : G502gat;
assign muxed225 = keyinput225 ? muxed254 : muxed213;
assign muxed226 = keyinput226 ? muxed203 : muxed257;
assign muxed227 = keyinput227 ? muxed359 : G330gat;
assign muxed228 = keyinput228 ? muxed164 : muxed359;
assign muxed229 = keyinput229 ? muxed204 : G853gat;
assign muxed230 = keyinput230 ? G625gat : muxed204;
assign muxed231 = keyinput231 ? muxed269 : G836gat;
assign muxed232 = keyinput232 ? muxed124 : G665gat;
assign muxed233 = keyinput233 ? muxed125 : G553gat;
assign muxed234 = keyinput234 ? muxed70 : muxed52;
assign muxed235 = keyinput235 ? G759gat : muxed70;
assign muxed236 = keyinput236 ? G624gat : G475gat;
assign muxed237 = keyinput237 ? G298gat : G624gat;
assign muxed238 = keyinput238 ? muxed31 : G585gat;
assign muxed239 = keyinput239 ? muxed271 : G761gat;
assign muxed240 = keyinput240 ? muxed382 : muxed271;
assign muxed241 = keyinput241 ? muxed273 : muxed204;
assign muxed242 = keyinput242 ? muxed211 : muxed276;
assign muxed243 = keyinput243 ? muxed57 : muxed276;
assign muxed244 = keyinput244 ? muxed384 : muxed57;
assign muxed245 = keyinput245 ? G490gat : G632gat;
assign muxed246 = keyinput246 ? G293gat : G490gat;
assign muxed247 = keyinput247 ? G751gat : muxed248;
assign muxed248 = keyinput248 ? G491gat : G712gat;
assign muxed249 = keyinput249 ? muxed223 : G379gat;
assign muxed250 = keyinput250 ? muxed224 : G477gat;
assign muxed251 = keyinput251 ? muxed290 : muxed164;
assign muxed252 = keyinput252 ? G376gat : muxed290;
assign muxed253 = keyinput253 ? muxed225 : muxed293;
assign muxed254 = keyinput254 ? G631gat : muxed14;
assign muxed255 = keyinput255 ? G507gat : G631gat;
assign muxed256 = keyinput256 ? muxed226 : G704gat;
assign muxed257 = keyinput257 ? G660gat : G324gat;
assign muxed258 = keyinput258 ? G552gat : G523gat;
assign muxed259 = keyinput259 ? G481gat : G552gat;
assign muxed260 = keyinput260 ? G530gat : muxed37;
assign muxed261 = keyinput261 ? muxed11 : G717gat;
assign muxed262 = keyinput262 ? G869gat : muxed11;
assign muxed263 = keyinput263 ? G842gat : G805gat;
assign muxed264 = keyinput264 ? muxed82 : G561gat;
assign muxed265 = keyinput265 ? G415gat : muxed82;
assign muxed266 = keyinput266 ? muxed17 : G586gat;
assign muxed267 = keyinput267 ? muxed49 : muxed64;
assign muxed268 = keyinput268 ? G781gat : G445gat;
assign muxed269 = keyinput269 ? G734gat : G781gat;
assign muxed270 = keyinput270 ? G51gat : muxed271;
assign muxed271 = keyinput271 ? muxed328 : muxed235;
assign muxed272 = keyinput272 ? muxed343 : G869gat;
assign muxed273 = keyinput273 ? muxed131 : G833gat;
assign muxed274 = keyinput274 ? muxed236 : muxed131;
assign muxed275 = keyinput275 ? muxed242 : G846gat;
assign muxed276 = keyinput276 ? G826gat : G722gat;
assign muxed277 = keyinput277 ? G808gat : muxed49;
assign muxed278 = keyinput278 ? G875gat : G808gat;
assign muxed279 = keyinput279 ? G802gat : muxed6;
assign muxed280 = keyinput280 ? muxed330 : G802gat;
assign muxed281 = keyinput281 ? muxed3 : muxed194;
assign muxed282 = keyinput282 ? muxed79 : muxed3;
assign muxed283 = keyinput283 ? muxed306 : G873gat;
assign muxed284 = keyinput284 ? muxed380 : muxed306;
assign muxed285 = keyinput285 ? muxed308 : muxed385;
assign muxed286 = keyinput286 ? muxed139 : G515gat;
assign muxed287 = keyinput287 ? muxed187 : muxed187;
assign muxed288 = keyinput288 ? muxed322 : G443gat;
assign muxed289 = keyinput289 ? muxed318 : muxed322;
assign muxed290 = keyinput290 ? muxed202 : G687gat;
assign muxed291 = keyinput291 ? muxed253 : muxed331;
assign muxed292 = keyinput292 ? muxed110 : muxed253;
assign muxed293 = keyinput293 ? G316gat : muxed142;
assign muxed294 = keyinput294 ? muxed150 : muxed346;
assign muxed295 = keyinput295 ? muxed327 : muxed349;
assign muxed296 = keyinput296 ? G814gat : muxed330;
assign muxed297 = keyinput297 ? muxed144 : G319gat;
assign muxed298 = keyinput298 ? muxed364 : muxed83;
assign muxed299 = keyinput299 ? muxed367 : muxed147;
assign muxed300 = keyinput300 ? muxed370 : G525gat;
assign muxed301 = keyinput301 ? muxed373 : G521gat;
assign muxed302 = keyinput302 ? muxed376 : G279gat;
assign muxed303 = keyinput303 ? muxed379 : G811gat;
assign muxed304 = keyinput304 ? muxed284 : muxed385;
assign muxed305 = keyinput305 ? G339gat : muxed284;
assign muxed306 = keyinput306 ? muxed169 : muxed70;
assign muxed307 = keyinput307 ? muxed285 : G743gat;
assign muxed308 = keyinput308 ? muxed186 : G764gat;
assign muxed309 = keyinput309 ? muxed62 : muxed186;
assign muxed310 = keyinput310 ? muxed88 : muxed179;
assign muxed311 = keyinput311 ? muxed262 : muxed88;
assign muxed312 = keyinput312 ? muxed170 : muxed286;
assign muxed313 = keyinput313 ? muxed323 : G516gat;
assign muxed314 = keyinput314 ? muxed252 : muxed323;
assign muxed315 = keyinput315 ? muxed96 : muxed316;
assign muxed316 = keyinput316 ? G460gat : G606gat;
assign muxed317 = keyinput317 ? G406gat : muxed188;
assign muxed318 = keyinput318 ? G303gat : G406gat;
assign muxed319 = keyinput319 ? G360gat : muxed9;
assign muxed320 = keyinput320 ? muxed289 : muxed231;
assign muxed321 = keyinput321 ? muxed34 : muxed289;
assign muxed322 = keyinput322 ? muxed314 : G512gat;
assign muxed323 = keyinput323 ? G847gat : G415gat;
assign muxed324 = keyinput324 ? muxed345 : muxed57;
assign muxed325 = keyinput325 ? G301gat : muxed345;
assign muxed326 = keyinput326 ? muxed347 : muxed334;
assign muxed327 = keyinput327 ? muxed92 : G498gat;
assign muxed328 = keyinput328 ? muxed210 : muxed92;
assign muxed329 = keyinput329 ? muxed296 : G752gat;
assign muxed330 = keyinput330 ? muxed291 : muxed374;
assign muxed331 = keyinput331 ? G533gat : G332gat;
assign muxed332 = keyinput332 ? muxed73 : G605gat;
assign muxed333 = keyinput333 ? muxed340 : muxed73;
assign muxed334 = keyinput334 ? G542gat : G338gat;
assign muxed335 = keyinput335 ? muxed74 : G745gat;
assign muxed336 = keyinput336 ? muxed282 : muxed74;
assign muxed337 = keyinput337 ? G437gat : G304gat;
assign muxed338 = keyinput338 ? muxed249 : muxed339;
assign muxed339 = keyinput339 ? muxed333 : G333gat;
assign muxed340 = keyinput340 ? G839gat : muxed5;
assign muxed341 = keyinput341 ? muxed245 : G839gat;
assign muxed342 = keyinput342 ? muxed221 : G857gat;
assign muxed343 = keyinput343 ? muxed241 : muxed221;
assign muxed344 = keyinput344 ? muxed325 : muxed12;
assign muxed345 = keyinput345 ? muxed294 : muxed169;
assign muxed346 = keyinput346 ? muxed326 : G871gat;
assign muxed347 = keyinput347 ? muxed295 : G764gat;
assign muxed348 = keyinput348 ? muxed119 : muxed295;
assign muxed349 = keyinput349 ? muxed45 : G651gat;
assign muxed350 = keyinput350 ? muxed215 : G415gat;
assign muxed351 = keyinput351 ? muxed133 : muxed198;
assign muxed352 = keyinput352 ? G295gat : muxed133;
assign muxed353 = keyinput353 ? muxed216 : muxed14;
assign muxed354 = keyinput354 ? G432gat : muxed216;
assign muxed355 = keyinput355 ? muxed220 : G298gat;
assign muxed356 = keyinput356 ? muxed86 : G502gat;
assign muxed357 = keyinput357 ? muxed100 : muxed86;
assign muxed358 = keyinput358 ? muxed228 : muxed6;
assign muxed359 = keyinput359 ? G569gat : G833gat;
assign muxed360 = keyinput360 ? muxed365 : muxed87;
assign muxed361 = keyinput361 ? muxed383 : muxed365;
assign muxed362 = keyinput362 ? G670gat : muxed363;
assign muxed363 = keyinput363 ? muxed298 : muxed29;
assign muxed364 = keyinput364 ? G793gat : G330gat;
assign muxed365 = keyinput365 ? G488gat : G793gat;
assign muxed366 = keyinput366 ? muxed299 : G498gat;
assign muxed367 = keyinput367 ? muxed145 : muxed328;
assign muxed368 = keyinput368 ? muxed134 : muxed145;
assign muxed369 = keyinput369 ? muxed300 : muxed157;
assign muxed370 = keyinput370 ? muxed112 : G285gat;
assign muxed371 = keyinput371 ? muxed10 : muxed112;
assign muxed372 = keyinput372 ? muxed301 : muxed3;
assign muxed373 = keyinput373 ? muxed178 : muxed164;
assign muxed374 = keyinput374 ? muxed268 : muxed178;
assign muxed375 = keyinput375 ? muxed302 : muxed19;
assign muxed376 = keyinput376 ? muxed160 : G628gat;
assign muxed377 = keyinput377 ? G732gat : muxed160;
assign muxed378 = keyinput378 ? muxed303 : G717gat;
assign muxed379 = keyinput379 ? muxed67 : G853gat;
assign muxed380 = keyinput380 ? G537gat : muxed67;
assign muxed381 = keyinput381 ? muxed361 : muxed144;
assign muxed382 = keyinput382 ? G848gat : muxed361;
assign muxed383 = keyinput383 ? muxed304 : muxed131;
assign muxed384 = keyinput384 ? muxed89 : muxed304;
assign muxed385 = keyinput385 ? muxed129 : muxed122;
assign muxed386 = keyinput386 ? G738gat : muxed96;
assign muxed387 = keyinput387 ? G856gat : G738gat;
endmodule
