`timescale 1ns / 1ps
// Verilog
// c880
// Ninputs 60
// Noutputs 26
// NtotalGates 383
// NAND4 13
// AND3 12
// NAND2 60
// NAND3 14
// AND2 105
// OR2 29
// NOT1 63
// NOR2 61
// BUFF1 26

module top (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
                  N865,N866,N874,N878,N879,N880,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
        keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
        keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
        keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
        keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
        keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
        keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
        keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
        keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
        keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
        keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
        keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
        keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
        keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
        keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
        keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
        keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
        keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
                  keyinput255,
        keyinput256, keyinput257, keyinput258, keyinput259, keyinput260,
        keyinput261, keyinput262, keyinput263, keyinput264, keyinput265,
        keyinput266, keyinput267, keyinput268, keyinput269, keyinput270,
        keyinput271, keyinput272, keyinput273, keyinput274, keyinput275,
        keyinput276, keyinput277, keyinput278, keyinput279, keyinput280,
        keyinput281, keyinput282, keyinput283, keyinput284, keyinput285,
        keyinput286, keyinput287, keyinput288, keyinput289, keyinput290,
        keyinput291, keyinput292, keyinput293, keyinput294, keyinput295,
        keyinput296, keyinput297, keyinput298, keyinput299, keyinput300,
        keyinput301, keyinput302, keyinput303, keyinput304, keyinput305,
        keyinput306, keyinput307, keyinput308, keyinput309, keyinput310,
        keyinput311, keyinput312, keyinput313, keyinput314, keyinput315,
        keyinput316, keyinput317, keyinput318, keyinput319, keyinput320,
        keyinput321, keyinput322, keyinput323, keyinput324, keyinput325,
        keyinput326, keyinput327, keyinput328, keyinput329, keyinput330,
        keyinput331, keyinput332, keyinput333, keyinput334, keyinput335,
        keyinput336, keyinput337, keyinput338, keyinput339, keyinput340,
        keyinput341, keyinput342, keyinput343, keyinput344, keyinput345,
        keyinput346, keyinput347, keyinput348, keyinput349, keyinput350,
        keyinput351, keyinput352, keyinput353, keyinput354, keyinput355,
        keyinput356, keyinput357, keyinput358, keyinput359, keyinput360,
        keyinput361, keyinput362, keyinput363, keyinput364, keyinput365,
        keyinput366, keyinput367, keyinput368, keyinput369, keyinput370,
                  keyinput371, keyinput372, keyinput373, keyinput374, keyinput375,
        keyinput376, keyinput377, keyinput378, keyinput379, keyinput380,
        keyinput381, keyinput382, keyinput383, keyinput384, keyinput385,
        keyinput386, keyinput387, keyinput388, keyinput389, keyinput390,
        keyinput391, keyinput392, keyinput393, keyinput394, keyinput395,
        keyinput396, keyinput397, keyinput398, keyinput399, keyinput400,
        keyinput401, keyinput402, keyinput403, keyinput404, keyinput405,
        keyinput406, keyinput407, keyinput408, keyinput409, keyinput410,
        keyinput411, keyinput412, keyinput413, keyinput414, keyinput415,
        keyinput416, keyinput417, keyinput418, keyinput419, keyinput420,
        keyinput421, keyinput422, keyinput423, keyinput424, keyinput425,
        keyinput426, keyinput427, keyinput428, keyinput429, keyinput430,
        keyinput431, keyinput432, keyinput433, keyinput434, keyinput435);

  input keyinput376, keyinput377, keyinput378, keyinput379, keyinput380;
  input keyinput381, keyinput382, keyinput383, keyinput384, keyinput385;
  input keyinput386, keyinput387, keyinput388, keyinput389, keyinput390;
  input keyinput391, keyinput392, keyinput393, keyinput394, keyinput395;
  input keyinput396, keyinput397, keyinput398, keyinput399, keyinput400;
  input keyinput401, keyinput402, keyinput403, keyinput404, keyinput405;
  input keyinput406, keyinput407, keyinput408, keyinput409, keyinput410;
  input keyinput411, keyinput412, keyinput413, keyinput414, keyinput415;
  input keyinput416, keyinput417, keyinput418, keyinput419, keyinput420;
  input keyinput421, keyinput422, keyinput423, keyinput424, keyinput425;
  input keyinput426, keyinput427, keyinput428, keyinput429, keyinput430;
  input keyinput431, keyinput432, keyinput433, keyinput434, keyinput435;


  input keyinput256, keyinput257, keyinput258, keyinput259, keyinput260;
  input keyinput261, keyinput262, keyinput263, keyinput264, keyinput265;
  input keyinput266, keyinput267, keyinput268, keyinput269, keyinput270;
  input keyinput271, keyinput272, keyinput273, keyinput274, keyinput275;
  input keyinput276, keyinput277, keyinput278, keyinput279, keyinput280;
  input keyinput281, keyinput282, keyinput283, keyinput284, keyinput285;
  input keyinput286, keyinput287, keyinput288, keyinput289, keyinput290;
  input keyinput291, keyinput292, keyinput293, keyinput294, keyinput295;
  input keyinput296, keyinput297, keyinput298, keyinput299, keyinput300;
  input keyinput301, keyinput302, keyinput303, keyinput304, keyinput305;
  input keyinput306, keyinput307, keyinput308, keyinput309, keyinput310;
  input keyinput311, keyinput312, keyinput313, keyinput314, keyinput315;
  input keyinput316, keyinput317, keyinput318, keyinput319, keyinput320;
  input keyinput321, keyinput322, keyinput323, keyinput324, keyinput325;
  input keyinput326, keyinput327, keyinput328, keyinput329, keyinput330;
  input keyinput331, keyinput332, keyinput333, keyinput334, keyinput335;
  input keyinput336, keyinput337, keyinput338, keyinput339, keyinput340;
  input keyinput341, keyinput342, keyinput343, keyinput344, keyinput345;
  input keyinput346, keyinput347, keyinput348, keyinput349, keyinput350;
  input keyinput351, keyinput352, keyinput353, keyinput354, keyinput355;
  input keyinput356, keyinput357, keyinput358, keyinput359, keyinput360;
  input keyinput361, keyinput362, keyinput363, keyinput364, keyinput365;
  input keyinput366, keyinput367, keyinput368, keyinput369, keyinput370;
  input keyinput371, keyinput372, keyinput373, keyinput374, keyinput375;

  wire KeyWire_0_1 , KeyWire_0_2, keyinput_Wire_1;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31, keyinput32, keyinput33, keyinput34;
  input keyinput35, keyinput36, keyinput37, keyinput38, keyinput39;
  input keyinput40, keyinput41, keyinput42, keyinput43, keyinput44;
  input keyinput45, keyinput46, keyinput47, keyinput48, keyinput49;
  input keyinput50, keyinput51, keyinput52, keyinput53, keyinput54;
  input keyinput55, keyinput56, keyinput57, keyinput58, keyinput59;
  input keyinput60, keyinput61, keyinput62, keyinput63, keyinput64;
  input keyinput65, keyinput66, keyinput67, keyinput68, keyinput69;
  input keyinput70, keyinput71, keyinput72, keyinput73, keyinput74;
  input keyinput75, keyinput76, keyinput77, keyinput78, keyinput79;
  input keyinput80, keyinput81, keyinput82, keyinput83, keyinput84;
  input keyinput85, keyinput86, keyinput87, keyinput88, keyinput89;
  input keyinput90, keyinput91, keyinput92, keyinput93, keyinput94;
  input keyinput95, keyinput96, keyinput97, keyinput98, keyinput99;
  input keyinput100, keyinput101, keyinput102, keyinput103, keyinput104;
  input keyinput105, keyinput106, keyinput107, keyinput108, keyinput109;
  input keyinput110, keyinput111, keyinput112, keyinput113, keyinput114;
  input keyinput115, keyinput116, keyinput117, keyinput118, keyinput119;
  input keyinput120, keyinput121, keyinput122, keyinput123, keyinput124;
  input keyinput125, keyinput126, keyinput127, keyinput128, keyinput129;
  input keyinput130, keyinput131, keyinput132, keyinput133, keyinput134;
  input keyinput135, keyinput136, keyinput137, keyinput138, keyinput139;
  input keyinput140, keyinput141, keyinput142, keyinput143, keyinput144;
  input keyinput145, keyinput146, keyinput147, keyinput148, keyinput149;
  input keyinput150, keyinput151, keyinput152, keyinput153, keyinput154;
  input keyinput155, keyinput156, keyinput157, keyinput158, keyinput159;
  input keyinput160, keyinput161, keyinput162, keyinput163, keyinput164;
  input keyinput165, keyinput166, keyinput167, keyinput168, keyinput169;
  input keyinput170, keyinput171, keyinput172, keyinput173, keyinput174;
  input keyinput175, keyinput176, keyinput177, keyinput178, keyinput179;
  input keyinput180, keyinput181, keyinput182, keyinput183, keyinput184;
  input keyinput185, keyinput186, keyinput187, keyinput188, keyinput189;
  input keyinput190, keyinput191, keyinput192, keyinput193, keyinput194;
  input keyinput195, keyinput196, keyinput197, keyinput198, keyinput199;
  input keyinput200, keyinput201, keyinput202, keyinput203, keyinput204;
  input keyinput205, keyinput206, keyinput207, keyinput208, keyinput209;
  input keyinput210, keyinput211, keyinput212, keyinput213, keyinput214;
  input keyinput215, keyinput216, keyinput217, keyinput218, keyinput219;
  input keyinput220, keyinput221, keyinput222, keyinput223, keyinput224;
  input keyinput225, keyinput226, keyinput227, keyinput228, keyinput229;
  input keyinput230, keyinput231, keyinput232, keyinput233, keyinput234;
  input keyinput235, keyinput236, keyinput237, keyinput238, keyinput239;
  input keyinput240, keyinput241, keyinput242, keyinput243, keyinput244;
  input keyinput245, keyinput246, keyinput247, keyinput248, keyinput249;
  input keyinput250, keyinput251, keyinput252, keyinput253, keyinput254;
  input keyinput255;

  wire [0:255] keyinput_Wire_0;
  wire [0:113] KeyNOTWire_0;

input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;

output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;

wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877;

nand NAND4_1 (N269, N1, N8, N13, N17);
nand NAND4_2 (N270, N1, N26, N13, N17);
and AND3_3 (N273, N29, N36, N42);
  and AND3_4 (keyinput_Wire_0[0], N1, N26, N51);
  xor keyGate_0_0(KeyNOTWire_0[0], keyinput0, keyinput_Wire_0[0]);
  not KeyNOTGate_0_0(N276, KeyNOTWire_0[0]);
  nand NAND4_5 (keyinput_Wire_0[1], N1, N8, N51, N17);
  xnor keyGate_0_1(KeyNOTWire_0[1], keyinput1, keyinput_Wire_0[1]);
  not KeyNOTGate_0_1(N279, KeyNOTWire_0[1]);
  nand NAND4_6 (keyinput_Wire_0[2], N1, N8, N13, N55);
  xor keyGate_0_2(KeyNOTWire_0[2], keyinput2, keyinput_Wire_0[2]);
  not KeyNOTGate_0_2(N280, KeyNOTWire_0[2]);
  nand NAND4_7 (keyinput_Wire_0[3], N59, N42, N68, N72);
  xor keyGate_0_3(KeyNOTWire_0[3], keyinput3, keyinput_Wire_0[3]);
  not KeyNOTGate_0_3(N284, KeyNOTWire_0[3]);
nand NAND2_8 (N285, N29, N68);
nand NAND3_9 (N286, N59, N68, N74);
  and AND3_10 (keyinput_Wire_0[4], N29, N75, N80);
  xor keyGate_0_4(N287, keyinput4, keyinput_Wire_0[4]);
and AND3_11 (N290, N29, N75, N42);
and AND3_12 (N291, N29, N36, N80);
and AND3_13 (N292, N29, N36, N42);
and AND3_14 (N293, N59, N75, N80);
  and AND3_15 (keyinput_Wire_0[5], N59, N75, N42);
  xnor keyGate_0_5(KeyNOTWire_0[4], keyinput5, keyinput_Wire_0[5]);
  not KeyNOTGate_0_4(N294, KeyNOTWire_0[4]);
and AND3_16 (N295, N59, N36, N80);
and AND3_17 (N296, N59, N36, N42);
and AND2_18 (N297, N85, N86);
or OR2_19 (N298, N87, N88);
nand NAND2_20 (N301, N91, N96);
or OR2_21 (N302, N91, N96);
nand NAND2_22 (N303, N101, N106);
or OR2_23 (N304, N101, N106);
nand NAND2_24 (N305, N111, N116);
or OR2_25 (N306, N111, N116);
nand NAND2_26 (N307, N121, N126);
or OR2_27 (N308, N121, N126);
and AND2_28 (N309, N8, N138);
  not NOT1_29 (keyinput_Wire_0[6], N268);
  xnor keyGate_0_6(KeyNOTWire_0[5], keyinput6, keyinput_Wire_0[6]);
  not KeyNOTGate_0_5(N310, KeyNOTWire_0[5]);
  and AND2_30 (keyinput_Wire_0[7], N51, N138);
  xor keyGate_0_7(N316, keyinput7, keyinput_Wire_0[7]);
  and AND2_31 (keyinput_Wire_0[8], N17, N138);
  xor keyGate_0_8(KeyNOTWire_0[6], keyinput8, keyinput_Wire_0[8]);
  not KeyNOTGate_0_6(N317, KeyNOTWire_0[6]);
  and AND2_32 (keyinput_Wire_0[9], N152, N138);
  xor keyGate_0_9(N318, keyinput9, keyinput_Wire_0[9]);
  nand NAND2_33 (keyinput_Wire_0[10], N59, N156);
  xnor keyGate_0_10(KeyNOTWire_0[7], keyinput10, keyinput_Wire_0[10]);
  not KeyNOTGate_0_7(N319, KeyNOTWire_0[7]);
  nor NOR2_34 (keyinput_Wire_0[11], N17, N42);
  xor keyGate_0_11(N322, keyinput11, keyinput_Wire_0[11]);
  and AND2_35 (keyinput_Wire_0[12], N17, N42);
  xor keyGate_0_12(N323, keyinput12, keyinput_Wire_0[12]);
nand NAND2_36 (N324, N159, N165);
or OR2_37 (N325, N159, N165);
nand NAND2_38 (N326, N171, N177);
or OR2_39 (N327, N171, N177);
nand NAND2_40 (N328, N183, N189);
or OR2_41 (N329, N183, N189);
nand NAND2_42 (N330, N195, N201);
or OR2_43 (N331, N195, N201);
and AND2_44 (N332, N210, N91);
and AND2_45 (N333, N210, N96);
and AND2_46 (N334, N210, N101);
and AND2_47 (N335, N210, N106);
and AND2_48 (N336, N210, N111);
and AND2_49 (N337, N255, N259);
and AND2_50 (N338, N210, N116);
and AND2_51 (N339, N255, N260);
and AND2_52 (N340, N210, N121);
and AND2_53 (N341, N255, N267);
not NOT1_54 (N342, N269);
not NOT1_55 (N343, N273);
or OR2_56 (N344, N270, N273);
  not NOT1_57 (keyinput_Wire_0[13], N276);
  xnor keyGate_0_13(N345, keyinput13, keyinput_Wire_0[13]);
not NOT1_58 (N346, N276);
  not NOT1_59 (keyinput_Wire_0[14], N279);
  xnor keyGate_0_14(N347, keyinput14, keyinput_Wire_0[14]);
  nor NOR2_60 (keyinput_Wire_0[15], N280, N284);
  xor keyGate_0_15(KeyNOTWire_0[8], keyinput15, keyinput_Wire_0[15]);
  not KeyNOTGate_0_8(N348, KeyNOTWire_0[8]);
or OR2_61 (N349, N280, N285);
or OR2_62 (N350, N280, N286);
not NOT1_63 (N351, N293);
  not NOT1_64 (keyinput_Wire_0[16], N294);
  xor keyGate_0_16(KeyNOTWire_0[9], keyinput16, keyinput_Wire_0[16]);
  not KeyNOTGate_0_9(N352, KeyNOTWire_0[9]);
not NOT1_65 (N353, N295);
not NOT1_66 (N354, N296);
nand NAND2_67 (N355, N89, N298);
and AND2_68 (N356, N90, N298);
nand NAND2_69 (N357, N301, N302);
nand NAND2_70 (N360, N303, N304);
nand NAND2_71 (N363, N305, N306);
nand NAND2_72 (N366, N307, N308);
  not NOT1_73 (keyinput_Wire_0[17], N310);
  xnor keyGate_0_17(N369, keyinput17, keyinput_Wire_0[17]);
  nor NOR2_74 (keyinput_Wire_0[18], N322, N323);
  xor keyGate_0_18(N375, keyinput18, keyinput_Wire_0[18]);
nand NAND2_75 (N376, N324, N325);
nand NAND2_76 (N379, N326, N327);
nand NAND2_77 (N382, N328, N329);
nand NAND2_78 (N385, N330, N331);
buf BUFF1_79 (N388, N290);
buf BUFF1_80 (N389, N291);
buf BUFF1_81 (N390, N292);
buf BUFF1_82 (N391, N297);
or OR2_83 (N392, N270, N343);
  not NOT1_84 (keyinput_Wire_0[19], N345);
  xnor keyGate_0_19(N393, keyinput19, keyinput_Wire_0[19]);
not NOT1_85 (N399, N346);
  and AND2_86 (keyinput_Wire_0[20], N348, N73);
  xor keyGate_0_20(KeyNOTWire_0[10], keyinput20, keyinput_Wire_0[20]);
  not KeyNOTGate_0_10(N400, KeyNOTWire_0[10]);
not NOT1_87 (N401, N349);
not NOT1_88 (N402, N350);
not NOT1_89 (N403, N355);
not NOT1_90 (N404, N357);
not NOT1_91 (N405, N360);
and AND2_92 (N406, N357, N360);
not NOT1_93 (N407, N363);
not NOT1_94 (N408, N366);
and AND2_95 (N409, N363, N366);
  nand NAND2_96 (keyinput_Wire_0[21], N347, N352);
  xnor keyGate_0_21(KeyNOTWire_0[11], keyinput21, keyinput_Wire_0[21]);
  not KeyNOTGate_0_11(N410, KeyNOTWire_0[11]);
not NOT1_97 (N411, N376);
not NOT1_98 (N412, N379);
and AND2_99 (N413, N376, N379);
not NOT1_100 (N414, N382);
not NOT1_101 (N415, N385);
and AND2_102 (N416, N382, N385);
and AND2_103 (N417, N210, N369);
buf BUFF1_104 (N418, N342);
buf BUFF1_105 (KeyWire_0_1, N344);
  xor flip_it (N419, KeyWire_0_1, KeyWire_0_2 );
buf BUFF1_106 (N420, N351);
buf BUFF1_107 (N421, N353);
buf BUFF1_108 (N422, N354);
buf BUFF1_109 (N423, N356);
  not NOT1_110 (keyinput_Wire_0[22], N400);
  xor keyGate_0_22(N424, keyinput22, keyinput_Wire_0[22]);
and AND2_111 (N425, N404, N405);
and AND2_112 (N426, N407, N408);
  and AND3_113 (keyinput_Wire_0[23], N319, N393, N55);
  xnor keyGate_0_23(N427, keyinput23, keyinput_Wire_0[23]);
  and AND3_114 (keyinput_Wire_0[24], N393, N17, N287);
  xnor keyGate_0_24(N432, keyinput24, keyinput_Wire_0[24]);
  nand NAND3_115 (keyinput_Wire_0[25], N393, N287, N55);
  xor keyGate_0_25(N437, keyinput25, keyinput_Wire_0[25]);
  nand NAND4_116 (keyinput_Wire_0[26], N375, N59, N156, N393);
  xor keyGate_0_26(KeyNOTWire_0[12], keyinput26, keyinput_Wire_0[26]);
  not KeyNOTGate_0_12(N442, KeyNOTWire_0[12]);
  nand NAND3_117 (keyinput_Wire_0[27], N393, N319, N17);
  xor keyGate_0_27(KeyNOTWire_0[13], keyinput27, keyinput_Wire_0[27]);
  not KeyNOTGate_0_13(N443, KeyNOTWire_0[13]);
and AND2_118 (N444, N411, N412);
and AND2_119 (N445, N414, N415);
buf BUFF1_120 (N446, N392);
buf BUFF1_121 (N447, N399);
buf BUFF1_122 (N448, N401);
buf BUFF1_123 (N449, N402);
buf BUFF1_124 (N450, N403);
  not NOT1_125 (keyinput_Wire_0[28], N424);
  xor keyGate_0_28(N451, keyinput28, keyinput_Wire_0[28]);
nor NOR2_126 (N460, N406, N425);
nor NOR2_127 (N463, N409, N426);
  nand NAND2_128 (keyinput_Wire_0[29], N442, N410);
  xnor keyGate_0_29(N466, keyinput29, keyinput_Wire_0[29]);
  and AND2_129 (keyinput_Wire_0[30], N143, N427);
  xnor keyGate_0_30(N475, keyinput30, keyinput_Wire_0[30]);
  and AND2_130 (keyinput_Wire_0[31], N310, N432);
  xor keyGate_0_31(N476, keyinput31, keyinput_Wire_0[31]);
  and AND2_131 (keyinput_Wire_0[32], N146, N427);
  xor keyGate_0_32(N477, keyinput32, keyinput_Wire_0[32]);
  and AND2_132 (keyinput_Wire_0[33], N310, N432);
  xor keyGate_0_33(N478, keyinput33, keyinput_Wire_0[33]);
  and AND2_133 (keyinput_Wire_0[34], N149, N427);
  xor keyGate_0_34(KeyNOTWire_0[14], keyinput34, keyinput_Wire_0[34]);
  not KeyNOTGate_0_14(N479, KeyNOTWire_0[14]);
  and AND2_134 (keyinput_Wire_0[35], N310, N432);
  xor keyGate_0_35(KeyNOTWire_0[15], keyinput35, keyinput_Wire_0[35]);
  not KeyNOTGate_0_15(N480, KeyNOTWire_0[15]);
  and AND2_135 (keyinput_Wire_0[36], N153, N427);
  xor keyGate_0_36(KeyNOTWire_0[16], keyinput36, keyinput_Wire_0[36]);
  not KeyNOTGate_0_16(N481, KeyNOTWire_0[16]);
  and AND2_136 (keyinput_Wire_0[37], N310, N432);
  xor keyGate_0_37(KeyNOTWire_0[17], keyinput37, keyinput_Wire_0[37]);
  not KeyNOTGate_0_17(N482, KeyNOTWire_0[17]);
  nand NAND2_137 (keyinput_Wire_0[38], N443, N1);
  xor keyGate_0_38(KeyNOTWire_0[18], keyinput38, keyinput_Wire_0[38]);
  not KeyNOTGate_0_18(N483, KeyNOTWire_0[18]);
  or OR2_138 (keyinput_Wire_0[39], N369, N437);
  xnor keyGate_0_39(N488, keyinput39, keyinput_Wire_0[39]);
  or OR2_139 (keyinput_Wire_0[40], N369, N437);
  xor keyGate_0_40(N489, keyinput40, keyinput_Wire_0[40]);
  or OR2_140 (keyinput_Wire_0[41], N369, N437);
  xor keyGate_0_41(KeyNOTWire_0[19], keyinput41, keyinput_Wire_0[41]);
  not KeyNOTGate_0_19(N490, KeyNOTWire_0[19]);
  or OR2_141 (keyinput_Wire_0[42], N369, N437);
  xor keyGate_0_42(N491, keyinput42, keyinput_Wire_0[42]);
nor NOR2_142 (N492, N413, N444);
nor NOR2_143 (N495, N416, N445);
nand NAND2_144 (N498, N130, N460);
or OR2_145 (N499, N130, N460);
nand NAND2_146 (N500, N463, N135);
or OR2_147 (N501, N463, N135);
  and AND2_148 (keyinput_Wire_0[43], N91, N466);
  xor keyGate_0_43(N502, keyinput43, keyinput_Wire_0[43]);
  nor NOR2_149 (keyinput_Wire_0[44], N475, N476);
  xnor keyGate_0_44(KeyNOTWire_0[20], keyinput44, keyinput_Wire_0[44]);
  not KeyNOTGate_0_20(N503, KeyNOTWire_0[20]);
  and AND2_150 (keyinput_Wire_0[45], N96, N466);
  xor keyGate_0_45(KeyNOTWire_0[21], keyinput45, keyinput_Wire_0[45]);
  not KeyNOTGate_0_21(N504, KeyNOTWire_0[21]);
  nor NOR2_151 (keyinput_Wire_0[46], N477, N478);
  xor keyGate_0_46(KeyNOTWire_0[22], keyinput46, keyinput_Wire_0[46]);
  not KeyNOTGate_0_22(N505, KeyNOTWire_0[22]);
  and AND2_152 (keyinput_Wire_0[47], N101, N466);
  xor keyGate_0_47(N506, keyinput47, keyinput_Wire_0[47]);
  nor NOR2_153 (keyinput_Wire_0[48], N479, N480);
  xor keyGate_0_48(N507, keyinput48, keyinput_Wire_0[48]);
  and AND2_154 (keyinput_Wire_0[49], N106, N466);
  xnor keyGate_0_49(N508, keyinput49, keyinput_Wire_0[49]);
  nor NOR2_155 (keyinput_Wire_0[50], N481, N482);
  xor keyGate_0_50(KeyNOTWire_0[23], keyinput50, keyinput_Wire_0[50]);
  not KeyNOTGate_0_23(N509, KeyNOTWire_0[23]);
  and AND2_156 (keyinput_Wire_0[51], N143, N483);
  xnor keyGate_0_51(N510, keyinput51, keyinput_Wire_0[51]);
  and AND2_157 (keyinput_Wire_0[52], N111, N466);
  xnor keyGate_0_52(KeyNOTWire_0[24], keyinput52, keyinput_Wire_0[52]);
  not KeyNOTGate_0_24(N511, KeyNOTWire_0[24]);
  and AND2_158 (keyinput_Wire_0[53], N146, N483);
  xnor keyGate_0_53(N512, keyinput53, keyinput_Wire_0[53]);
  and AND2_159 (keyinput_Wire_0[54], N116, N466);
  xor keyGate_0_54(KeyNOTWire_0[25], keyinput54, keyinput_Wire_0[54]);
  not KeyNOTGate_0_25(N513, KeyNOTWire_0[25]);
  and AND2_160 (keyinput_Wire_0[55], N149, N483);
  xor keyGate_0_55(KeyNOTWire_0[26], keyinput55, keyinput_Wire_0[55]);
  not KeyNOTGate_0_26(N514, KeyNOTWire_0[26]);
  and AND2_161 (keyinput_Wire_0[56], N121, N466);
  xnor keyGate_0_56(N515, keyinput56, keyinput_Wire_0[56]);
  and AND2_162 (keyinput_Wire_0[57], N153, N483);
  xnor keyGate_0_57(KeyNOTWire_0[27], keyinput57, keyinput_Wire_0[57]);
  not KeyNOTGate_0_27(N516, KeyNOTWire_0[27]);
  and AND2_163 (keyinput_Wire_0[58], N126, N466);
  xnor keyGate_0_58(N517, keyinput58, keyinput_Wire_0[58]);
nand NAND2_164 (N518, N130, N492);
or OR2_165 (N519, N130, N492);
nand NAND2_166 (N520, N495, N207);
or OR2_167 (N521, N495, N207);
and AND2_168 (N522, N451, N159);
and AND2_169 (N523, N451, N165);
and AND2_170 (N524, N451, N171);
and AND2_171 (N525, N451, N177);
and AND2_172 (N526, N451, N183);
nand NAND2_173 (N527, N451, N189);
nand NAND2_174 (N528, N451, N195);
nand NAND2_175 (N529, N451, N201);
  nand NAND2_176 (keyinput_Wire_0[59], N498, N499);
  xnor keyGate_0_59(N530, keyinput59, keyinput_Wire_0[59]);
  nand NAND2_177 (keyinput_Wire_0[60], N500, N501);
  xor keyGate_0_60(N533, keyinput60, keyinput_Wire_0[60]);
  nor NOR2_178 (keyinput_Wire_0[61], N309, N502);
  xor keyGate_0_61(N536, keyinput61, keyinput_Wire_0[61]);
  nor NOR2_179 (keyinput_Wire_0[62], N316, N504);
  xnor keyGate_0_62(KeyNOTWire_0[28], keyinput62, keyinput_Wire_0[62]);
  not KeyNOTGate_0_28(N537, KeyNOTWire_0[28]);
  nor NOR2_180 (keyinput_Wire_0[63], N317, N506);
  xor keyGate_0_63(N538, keyinput63, keyinput_Wire_0[63]);
  nor NOR2_181 (keyinput_Wire_0[64], N318, N508);
  xnor keyGate_0_64(N539, keyinput64, keyinput_Wire_0[64]);
  nor NOR2_182 (keyinput_Wire_0[65], N510, N511);
  xor keyGate_0_65(N540, keyinput65, keyinput_Wire_0[65]);
  nor NOR2_183 (keyinput_Wire_0[66], N512, N513);
  xor keyGate_0_66(KeyNOTWire_0[29], keyinput66, keyinput_Wire_0[66]);
  not KeyNOTGate_0_29(N541, KeyNOTWire_0[29]);
  nor NOR2_184 (keyinput_Wire_0[67], N514, N515);
  xnor keyGate_0_67(N542, keyinput67, keyinput_Wire_0[67]);
  nor NOR2_185 (keyinput_Wire_0[68], N516, N517);
  xor keyGate_0_68(KeyNOTWire_0[30], keyinput68, keyinput_Wire_0[68]);
  not KeyNOTGate_0_30(N543, KeyNOTWire_0[30]);
  nand NAND2_186 (keyinput_Wire_0[69], N518, N519);
  xor keyGate_0_69(KeyNOTWire_0[31], keyinput69, keyinput_Wire_0[69]);
  not KeyNOTGate_0_31(N544, KeyNOTWire_0[31]);
  nand NAND2_187 (keyinput_Wire_0[70], N520, N521);
  xnor keyGate_0_70(KeyNOTWire_0[32], keyinput70, keyinput_Wire_0[70]);
  not KeyNOTGate_0_32(N547, KeyNOTWire_0[32]);
  not NOT1_188 (keyinput_Wire_0[71], N530);
  xor keyGate_0_71(N550, keyinput71, keyinput_Wire_0[71]);
  not NOT1_189 (keyinput_Wire_0[72], N533);
  xnor keyGate_0_72(N551, keyinput72, keyinput_Wire_0[72]);
  and AND2_190 (keyinput_Wire_0[73], N530, N533);
  xnor keyGate_0_73(N552, keyinput73, keyinput_Wire_0[73]);
  nand NAND2_191 (keyinput_Wire_0[74], N536, N503);
  xnor keyGate_0_74(N553, keyinput74, keyinput_Wire_0[74]);
  nand NAND2_192 (keyinput_Wire_0[75], N537, N505);
  xnor keyGate_0_75(N557, keyinput75, keyinput_Wire_0[75]);
  nand NAND2_193 (keyinput_Wire_0[76], N538, N507);
  xnor keyGate_0_76(N561, keyinput76, keyinput_Wire_0[76]);
  nand NAND2_194 (keyinput_Wire_0[77], N539, N509);
  xor keyGate_0_77(N565, keyinput77, keyinput_Wire_0[77]);
  nand NAND2_195 (keyinput_Wire_0[78], N488, N540);
  xnor keyGate_0_78(N569, keyinput78, keyinput_Wire_0[78]);
  nand NAND2_196 (keyinput_Wire_0[79], N489, N541);
  xnor keyGate_0_79(N573, keyinput79, keyinput_Wire_0[79]);
  nand NAND2_197 (keyinput_Wire_0[80], N490, N542);
  xnor keyGate_0_80(N577, keyinput80, keyinput_Wire_0[80]);
  nand NAND2_198 (keyinput_Wire_0[81], N491, N543);
  xnor keyGate_0_81(N581, keyinput81, keyinput_Wire_0[81]);
  not NOT1_199 (keyinput_Wire_0[82], N544);
  xnor keyGate_0_82(N585, keyinput82, keyinput_Wire_0[82]);
  not NOT1_200 (keyinput_Wire_0[83], N547);
  xnor keyGate_0_83(KeyNOTWire_0[33], keyinput83, keyinput_Wire_0[83]);
  not KeyNOTGate_0_33(N586, KeyNOTWire_0[33]);
  and AND2_201 (keyinput_Wire_0[84], N544, N547);
  xor keyGate_0_84(KeyNOTWire_0[34], keyinput84, keyinput_Wire_0[84]);
  not KeyNOTGate_0_34(N587, KeyNOTWire_0[34]);
  and AND2_202 (keyinput_Wire_0[85], N550, N551);
  xor keyGate_0_85(N588, keyinput85, keyinput_Wire_0[85]);
  and AND2_203 (keyinput_Wire_0[86], N585, N586);
  xnor keyGate_0_86(KeyNOTWire_0[35], keyinput86, keyinput_Wire_0[86]);
  not KeyNOTGate_0_35(N589, KeyNOTWire_0[35]);
  nand NAND2_204 (keyinput_Wire_0[87], N553, N159);
  xnor keyGate_0_87(N590, keyinput87, keyinput_Wire_0[87]);
  or OR2_205 (keyinput_Wire_0[88], N553, N159);
  xor keyGate_0_88(N593, keyinput88, keyinput_Wire_0[88]);
  and AND2_206 (keyinput_Wire_0[89], N246, N553);
  xor keyGate_0_89(N596, keyinput89, keyinput_Wire_0[89]);
  nand NAND2_207 (keyinput_Wire_0[90], N557, N165);
  xnor keyGate_0_90(KeyNOTWire_0[36], keyinput90, keyinput_Wire_0[90]);
  not KeyNOTGate_0_36(N597, KeyNOTWire_0[36]);
  or OR2_208 (keyinput_Wire_0[91], N557, N165);
  xor keyGate_0_91(N600, keyinput91, keyinput_Wire_0[91]);
  and AND2_209 (keyinput_Wire_0[92], N246, N557);
  xnor keyGate_0_92(KeyNOTWire_0[37], keyinput92, keyinput_Wire_0[92]);
  not KeyNOTGate_0_37(N605, KeyNOTWire_0[37]);
  nand NAND2_210 (keyinput_Wire_0[93], N561, N171);
  xor keyGate_0_93(N606, keyinput93, keyinput_Wire_0[93]);
  or OR2_211 (keyinput_Wire_0[94], N561, N171);
  xor keyGate_0_94(KeyNOTWire_0[38], keyinput94, keyinput_Wire_0[94]);
  not KeyNOTGate_0_38(N609, KeyNOTWire_0[38]);
  and AND2_212 (keyinput_Wire_0[95], N246, N561);
  xor keyGate_0_95(N615, keyinput95, keyinput_Wire_0[95]);
  nand NAND2_213 (keyinput_Wire_0[96], N565, N177);
  xnor keyGate_0_96(KeyNOTWire_0[39], keyinput96, keyinput_Wire_0[96]);
  not KeyNOTGate_0_39(N616, KeyNOTWire_0[39]);
  or OR2_214 (keyinput_Wire_0[97], N565, N177);
  xor keyGate_0_97(KeyNOTWire_0[40], keyinput97, keyinput_Wire_0[97]);
  not KeyNOTGate_0_40(N619, KeyNOTWire_0[40]);
  and AND2_215 (keyinput_Wire_0[98], N246, N565);
  xnor keyGate_0_98(N624, keyinput98, keyinput_Wire_0[98]);
  nand NAND2_216 (keyinput_Wire_0[99], N569, N183);
  xnor keyGate_0_99(N625, keyinput99, keyinput_Wire_0[99]);
  or OR2_217 (keyinput_Wire_0[100], N569, N183);
  xnor keyGate_0_100(N628, keyinput100, keyinput_Wire_0[100]);
  and AND2_218 (keyinput_Wire_0[101], N246, N569);
  xnor keyGate_0_101(KeyNOTWire_0[41], keyinput101, keyinput_Wire_0[101]);
  not KeyNOTGate_0_41(N631, KeyNOTWire_0[41]);
  nand NAND2_219 (keyinput_Wire_0[102], N573, N189);
  xor keyGate_0_102(KeyNOTWire_0[42], keyinput102, keyinput_Wire_0[102]);
  not KeyNOTGate_0_42(N632, KeyNOTWire_0[42]);
  or OR2_220 (keyinput_Wire_0[103], N573, N189);
  xnor keyGate_0_103(N635, keyinput103, keyinput_Wire_0[103]);
  and AND2_221 (keyinput_Wire_0[104], N246, N573);
  xor keyGate_0_104(N640, keyinput104, keyinput_Wire_0[104]);
  nand NAND2_222 (keyinput_Wire_0[105], N577, N195);
  xor keyGate_0_105(KeyNOTWire_0[43], keyinput105, keyinput_Wire_0[105]);
  not KeyNOTGate_0_43(N641, KeyNOTWire_0[43]);
  or OR2_223 (keyinput_Wire_0[106], N577, N195);
  xnor keyGate_0_106(N644, keyinput106, keyinput_Wire_0[106]);
  and AND2_224 (keyinput_Wire_0[107], N246, N577);
  xnor keyGate_0_107(N650, keyinput107, keyinput_Wire_0[107]);
  nand NAND2_225 (keyinput_Wire_0[108], N581, N201);
  xor keyGate_0_108(N651, keyinput108, keyinput_Wire_0[108]);
  or OR2_226 (keyinput_Wire_0[109], N581, N201);
  xnor keyGate_0_109(N654, keyinput109, keyinput_Wire_0[109]);
  and AND2_227 (keyinput_Wire_0[110], N246, N581);
  xor keyGate_0_110(KeyNOTWire_0[44], keyinput110, keyinput_Wire_0[110]);
  not KeyNOTGate_0_44(N659, KeyNOTWire_0[44]);
  nor NOR2_228 (keyinput_Wire_0[111], N552, N588);
  xor keyGate_0_111(KeyNOTWire_0[45], keyinput111, keyinput_Wire_0[111]);
  not KeyNOTGate_0_45(N660, KeyNOTWire_0[45]);
  nor NOR2_229 (keyinput_Wire_0[112], N587, N589);
  xnor keyGate_0_112(N661, keyinput112, keyinput_Wire_0[112]);
  not NOT1_230 (keyinput_Wire_0[113], N590);
  xnor keyGate_0_113(N662, keyinput113, keyinput_Wire_0[113]);
  and AND2_231 (keyinput_Wire_0[114], N593, N590);
  xor keyGate_0_114(KeyNOTWire_0[46], keyinput114, keyinput_Wire_0[114]);
  not KeyNOTGate_0_46(N665, KeyNOTWire_0[46]);
  nor NOR2_232 (keyinput_Wire_0[115], N596, N522);
  xnor keyGate_0_115(KeyNOTWire_0[47], keyinput115, keyinput_Wire_0[115]);
  not KeyNOTGate_0_47(N669, KeyNOTWire_0[47]);
  not NOT1_233 (keyinput_Wire_0[116], N597);
  xnor keyGate_0_116(N670, keyinput116, keyinput_Wire_0[116]);
  and AND2_234 (keyinput_Wire_0[117], N600, N597);
  xor keyGate_0_117(N673, keyinput117, keyinput_Wire_0[117]);
  nor NOR2_235 (keyinput_Wire_0[118], N605, N523);
  xnor keyGate_0_118(KeyNOTWire_0[48], keyinput118, keyinput_Wire_0[118]);
  not KeyNOTGate_0_48(N677, KeyNOTWire_0[48]);
  not NOT1_236 (keyinput_Wire_0[119], N606);
  xor keyGate_0_119(KeyNOTWire_0[49], keyinput119, keyinput_Wire_0[119]);
  not KeyNOTGate_0_49(N678, KeyNOTWire_0[49]);
  and AND2_237 (keyinput_Wire_0[120], N609, N606);
  xnor keyGate_0_120(N682, keyinput120, keyinput_Wire_0[120]);
  nor NOR2_238 (keyinput_Wire_0[121], N615, N524);
  xor keyGate_0_121(N686, keyinput121, keyinput_Wire_0[121]);
  not NOT1_239 (keyinput_Wire_0[122], N616);
  xor keyGate_0_122(N687, keyinput122, keyinput_Wire_0[122]);
  and AND2_240 (keyinput_Wire_0[123], N619, N616);
  xnor keyGate_0_123(N692, keyinput123, keyinput_Wire_0[123]);
  nor NOR2_241 (keyinput_Wire_0[124], N624, N525);
  xnor keyGate_0_124(KeyNOTWire_0[50], keyinput124, keyinput_Wire_0[124]);
  not KeyNOTGate_0_50(N696, KeyNOTWire_0[50]);
  not NOT1_242 (keyinput_Wire_0[125], N625);
  xor keyGate_0_125(KeyNOTWire_0[51], keyinput125, keyinput_Wire_0[125]);
  not KeyNOTGate_0_51(N697, KeyNOTWire_0[51]);
  and AND2_243 (keyinput_Wire_0[126], N628, N625);
  xnor keyGate_0_126(KeyNOTWire_0[52], keyinput126, keyinput_Wire_0[126]);
  not KeyNOTGate_0_52(N700, KeyNOTWire_0[52]);
  nor NOR2_244 (keyinput_Wire_0[127], N631, N526);
  xnor keyGate_0_127(KeyNOTWire_0[53], keyinput127, keyinput_Wire_0[127]);
  not KeyNOTGate_0_53(N704, KeyNOTWire_0[53]);
  not NOT1_245 (keyinput_Wire_0[128], N632);
  xor keyGate_0_128(KeyNOTWire_0[54], keyinput128, keyinput_Wire_0[128]);
  not KeyNOTGate_0_54(N705, KeyNOTWire_0[54]);
  and AND2_246 (keyinput_Wire_0[129], N635, N632);
  xor keyGate_0_129(N708, keyinput129, keyinput_Wire_0[129]);
  nor NOR2_247 (keyinput_Wire_0[130], N337, N640);
  xor keyGate_0_130(N712, keyinput130, keyinput_Wire_0[130]);
  not NOT1_248 (keyinput_Wire_0[131], N641);
  xnor keyGate_0_131(N713, keyinput131, keyinput_Wire_0[131]);
  and AND2_249 (keyinput_Wire_0[132], N644, N641);
  xnor keyGate_0_132(KeyNOTWire_0[55], keyinput132, keyinput_Wire_0[132]);
  not KeyNOTGate_0_55(N717, KeyNOTWire_0[55]);
  nor NOR2_250 (keyinput_Wire_0[133], N339, N650);
  xnor keyGate_0_133(N721, keyinput133, keyinput_Wire_0[133]);
  not NOT1_251 (keyinput_Wire_0[134], N651);
  xnor keyGate_0_134(N722, keyinput134, keyinput_Wire_0[134]);
  and AND2_252 (keyinput_Wire_0[135], N654, N651);
  xor keyGate_0_135(N727, keyinput135, keyinput_Wire_0[135]);
  nor NOR2_253 (keyinput_Wire_0[136], N341, N659);
  xor keyGate_0_136(KeyNOTWire_0[56], keyinput136, keyinput_Wire_0[136]);
  not KeyNOTGate_0_56(N731, KeyNOTWire_0[56]);
  nand NAND2_254 (keyinput_Wire_0[137], N654, N261);
  xnor keyGate_0_137(KeyNOTWire_0[57], keyinput137, keyinput_Wire_0[137]);
  not KeyNOTGate_0_57(N732, KeyNOTWire_0[57]);
  nand NAND3_255 (keyinput_Wire_0[138], N644, N654, N261);
  xnor keyGate_0_138(N733, keyinput138, keyinput_Wire_0[138]);
  nand NAND4_256 (keyinput_Wire_0[139], N635, N644, N654, N261);
  xor keyGate_0_139(KeyNOTWire_0[58], keyinput139, keyinput_Wire_0[139]);
  not KeyNOTGate_0_58(N734, KeyNOTWire_0[58]);
  not NOT1_257 (keyinput_Wire_0[140], N662);
  xor keyGate_0_140(KeyNOTWire_0[59], keyinput140, keyinput_Wire_0[140]);
  not KeyNOTGate_0_59(N735, KeyNOTWire_0[59]);
  and AND2_258 (keyinput_Wire_0[141], N228, N665);
  xor keyGate_0_141(KeyNOTWire_0[60], keyinput141, keyinput_Wire_0[141]);
  not KeyNOTGate_0_60(N736, KeyNOTWire_0[60]);
  and AND2_259 (keyinput_Wire_0[142], N237, N662);
  xor keyGate_0_142(KeyNOTWire_0[61], keyinput142, keyinput_Wire_0[142]);
  not KeyNOTGate_0_61(N737, KeyNOTWire_0[61]);
  not NOT1_260 (keyinput_Wire_0[143], N670);
  xnor keyGate_0_143(N738, keyinput143, keyinput_Wire_0[143]);
  and AND2_261 (keyinput_Wire_0[144], N228, N673);
  xor keyGate_0_144(N739, keyinput144, keyinput_Wire_0[144]);
  and AND2_262 (keyinput_Wire_0[145], N237, N670);
  xor keyGate_0_145(KeyNOTWire_0[62], keyinput145, keyinput_Wire_0[145]);
  not KeyNOTGate_0_62(N740, KeyNOTWire_0[62]);
  not NOT1_263 (keyinput_Wire_0[146], N678);
  xor keyGate_0_146(KeyNOTWire_0[63], keyinput146, keyinput_Wire_0[146]);
  not KeyNOTGate_0_63(N741, KeyNOTWire_0[63]);
  and AND2_264 (keyinput_Wire_0[147], N228, N682);
  xnor keyGate_0_147(N742, keyinput147, keyinput_Wire_0[147]);
  and AND2_265 (keyinput_Wire_0[148], N237, N678);
  xnor keyGate_0_148(KeyNOTWire_0[64], keyinput148, keyinput_Wire_0[148]);
  not KeyNOTGate_0_64(N743, KeyNOTWire_0[64]);
  not NOT1_266 (keyinput_Wire_0[149], N687);
  xnor keyGate_0_149(KeyNOTWire_0[65], keyinput149, keyinput_Wire_0[149]);
  not KeyNOTGate_0_65(N744, KeyNOTWire_0[65]);
  and AND2_267 (keyinput_Wire_0[150], N228, N692);
  xor keyGate_0_150(N745, keyinput150, keyinput_Wire_0[150]);
  and AND2_268 (keyinput_Wire_0[151], N237, N687);
  xor keyGate_0_151(N746, keyinput151, keyinput_Wire_0[151]);
  not NOT1_269 (keyinput_Wire_0[152], N697);
  xor keyGate_0_152(N747, keyinput152, keyinput_Wire_0[152]);
  and AND2_270 (keyinput_Wire_0[153], N228, N700);
  xnor keyGate_0_153(N748, keyinput153, keyinput_Wire_0[153]);
  and AND2_271 (keyinput_Wire_0[154], N237, N697);
  xor keyGate_0_154(N749, keyinput154, keyinput_Wire_0[154]);
  not NOT1_272 (keyinput_Wire_0[155], N705);
  xor keyGate_0_155(N750, keyinput155, keyinput_Wire_0[155]);
  and AND2_273 (keyinput_Wire_0[156], N228, N708);
  xor keyGate_0_156(N751, keyinput156, keyinput_Wire_0[156]);
  and AND2_274 (keyinput_Wire_0[157], N237, N705);
  xnor keyGate_0_157(KeyNOTWire_0[66], keyinput157, keyinput_Wire_0[157]);
  not KeyNOTGate_0_66(N752, KeyNOTWire_0[66]);
  not NOT1_275 (keyinput_Wire_0[158], N713);
  xnor keyGate_0_158(N753, keyinput158, keyinput_Wire_0[158]);
  and AND2_276 (keyinput_Wire_0[159], N228, N717);
  xnor keyGate_0_159(KeyNOTWire_0[67], keyinput159, keyinput_Wire_0[159]);
  not KeyNOTGate_0_67(N754, KeyNOTWire_0[67]);
  and AND2_277 (keyinput_Wire_0[160], N237, N713);
  xor keyGate_0_160(N755, keyinput160, keyinput_Wire_0[160]);
  not NOT1_278 (keyinput_Wire_0[161], N722);
  xnor keyGate_0_161(N756, keyinput161, keyinput_Wire_0[161]);
  nor NOR2_279 (keyinput_Wire_0[162], N727, N261);
  xor keyGate_0_162(KeyNOTWire_0[68], keyinput162, keyinput_Wire_0[162]);
  not KeyNOTGate_0_68(N757, KeyNOTWire_0[68]);
  and AND2_280 (keyinput_Wire_0[163], N727, N261);
  xor keyGate_0_163(KeyNOTWire_0[69], keyinput163, keyinput_Wire_0[163]);
  not KeyNOTGate_0_69(N758, KeyNOTWire_0[69]);
  and AND2_281 (keyinput_Wire_0[164], N228, N727);
  xnor keyGate_0_164(KeyNOTWire_0[70], keyinput164, keyinput_Wire_0[164]);
  not KeyNOTGate_0_70(N759, KeyNOTWire_0[70]);
  and AND2_282 (keyinput_Wire_0[165], N237, N722);
  xor keyGate_0_165(KeyNOTWire_0[71], keyinput165, keyinput_Wire_0[165]);
  not KeyNOTGate_0_71(N760, KeyNOTWire_0[71]);
  nand NAND2_283 (keyinput_Wire_0[166], N644, N722);
  xor keyGate_0_166(KeyNOTWire_0[72], keyinput166, keyinput_Wire_0[166]);
  not KeyNOTGate_0_72(N761, KeyNOTWire_0[72]);
  nand NAND2_284 (keyinput_Wire_0[167], N635, N713);
  xor keyGate_0_167(N762, keyinput167, keyinput_Wire_0[167]);
  nand NAND3_285 (keyinput_Wire_0[168], N635, N644, N722);
  xor keyGate_0_168(KeyNOTWire_0[73], keyinput168, keyinput_Wire_0[168]);
  not KeyNOTGate_0_73(N763, KeyNOTWire_0[73]);
  nand NAND2_286 (keyinput_Wire_0[169], N609, N687);
  xor keyGate_0_169(KeyNOTWire_0[74], keyinput169, keyinput_Wire_0[169]);
  not KeyNOTGate_0_74(N764, KeyNOTWire_0[74]);
  nand NAND2_287 (keyinput_Wire_0[170], N600, N678);
  xnor keyGate_0_170(KeyNOTWire_0[75], keyinput170, keyinput_Wire_0[170]);
  not KeyNOTGate_0_75(N765, KeyNOTWire_0[75]);
  nand NAND3_288 (keyinput_Wire_0[171], N600, N609, N687);
  xnor keyGate_0_171(N766, keyinput171, keyinput_Wire_0[171]);
buf BUFF1_289 (N767, N660);
buf BUFF1_290 (N768, N661);
  nor NOR2_291 (keyinput_Wire_0[172], N736, N737);
  xnor keyGate_0_172(KeyNOTWire_0[76], keyinput172, keyinput_Wire_0[172]);
  not KeyNOTGate_0_76(N769, KeyNOTWire_0[76]);
  nor NOR2_292 (keyinput_Wire_0[173], N739, N740);
  xor keyGate_0_173(KeyNOTWire_0[77], keyinput173, keyinput_Wire_0[173]);
  not KeyNOTGate_0_77(N770, KeyNOTWire_0[77]);
  nor NOR2_293 (keyinput_Wire_0[174], N742, N743);
  xor keyGate_0_174(N771, keyinput174, keyinput_Wire_0[174]);
  nor NOR2_294 (keyinput_Wire_0[175], N745, N746);
  xnor keyGate_0_175(N772, keyinput175, keyinput_Wire_0[175]);
  nand NAND4_295 (keyinput_Wire_0[176], N750, N762, N763, N734);
  xor keyGate_0_176(N773, keyinput176, keyinput_Wire_0[176]);
  nor NOR2_296 (keyinput_Wire_0[177], N748, N749);
  xnor keyGate_0_177(N777, keyinput177, keyinput_Wire_0[177]);
  nand NAND3_297 (keyinput_Wire_0[178], N753, N761, N733);
  xor keyGate_0_178(KeyNOTWire_0[78], keyinput178, keyinput_Wire_0[178]);
  not KeyNOTGate_0_78(N778, KeyNOTWire_0[78]);
  nor NOR2_298 (keyinput_Wire_0[179], N751, N752);
  xnor keyGate_0_179(N781, keyinput179, keyinput_Wire_0[179]);
  nand NAND2_299 (keyinput_Wire_0[180], N756, N732);
  xor keyGate_0_180(N782, keyinput180, keyinput_Wire_0[180]);
  nor NOR2_300 (keyinput_Wire_0[181], N754, N755);
  xnor keyGate_0_181(N785, keyinput181, keyinput_Wire_0[181]);
  nor NOR2_301 (keyinput_Wire_0[182], N757, N758);
  xnor keyGate_0_182(KeyNOTWire_0[79], keyinput182, keyinput_Wire_0[182]);
  not KeyNOTGate_0_79(N786, KeyNOTWire_0[79]);
  nor NOR2_302 (keyinput_Wire_0[183], N759, N760);
  xnor keyGate_0_183(N787, keyinput183, keyinput_Wire_0[183]);
  nor NOR2_303 (keyinput_Wire_0[184], N700, N773);
  xnor keyGate_0_184(KeyNOTWire_0[80], keyinput184, keyinput_Wire_0[184]);
  not KeyNOTGate_0_80(N788, KeyNOTWire_0[80]);
  and AND2_304 (keyinput_Wire_0[185], N700, N773);
  xor keyGate_0_185(N789, keyinput185, keyinput_Wire_0[185]);
  nor NOR2_305 (keyinput_Wire_0[186], N708, N778);
  xor keyGate_0_186(KeyNOTWire_0[81], keyinput186, keyinput_Wire_0[186]);
  not KeyNOTGate_0_81(N790, KeyNOTWire_0[81]);
  and AND2_306 (keyinput_Wire_0[187], N708, N778);
  xnor keyGate_0_187(N791, keyinput187, keyinput_Wire_0[187]);
  nor NOR2_307 (keyinput_Wire_0[188], N717, N782);
  xor keyGate_0_188(KeyNOTWire_0[82], keyinput188, keyinput_Wire_0[188]);
  not KeyNOTGate_0_82(N792, KeyNOTWire_0[82]);
  and AND2_308 (keyinput_Wire_0[189], N717, N782);
  xor keyGate_0_189(N793, keyinput189, keyinput_Wire_0[189]);
  and AND2_309 (keyinput_Wire_0[190], N219, N786);
  xnor keyGate_0_190(N794, keyinput190, keyinput_Wire_0[190]);
  nand NAND2_310 (keyinput_Wire_0[191], N628, N773);
  xor keyGate_0_191(N795, keyinput191, keyinput_Wire_0[191]);
  nand NAND2_311 (keyinput_Wire_0[192], N795, N747);
  xor keyGate_0_192(KeyNOTWire_0[83], keyinput192, keyinput_Wire_0[192]);
  not KeyNOTGate_0_83(N796, KeyNOTWire_0[83]);
  nor NOR2_312 (keyinput_Wire_0[193], N788, N789);
  xor keyGate_0_193(KeyNOTWire_0[84], keyinput193, keyinput_Wire_0[193]);
  not KeyNOTGate_0_84(N802, KeyNOTWire_0[84]);
  nor NOR2_313 (keyinput_Wire_0[194], N790, N791);
  xnor keyGate_0_194(KeyNOTWire_0[85], keyinput194, keyinput_Wire_0[194]);
  not KeyNOTGate_0_85(N803, KeyNOTWire_0[85]);
  nor NOR2_314 (keyinput_Wire_0[195], N792, N793);
  xor keyGate_0_195(N804, keyinput195, keyinput_Wire_0[195]);
  nor NOR2_315 (keyinput_Wire_0[196], N340, N794);
  xnor keyGate_0_196(N805, keyinput196, keyinput_Wire_0[196]);
  nor NOR2_316 (keyinput_Wire_0[197], N692, N796);
  xor keyGate_0_197(KeyNOTWire_0[86], keyinput197, keyinput_Wire_0[197]);
  not KeyNOTGate_0_86(N806, KeyNOTWire_0[86]);
  and AND2_317 (keyinput_Wire_0[198], N692, N796);
  xor keyGate_0_198(KeyNOTWire_0[87], keyinput198, keyinput_Wire_0[198]);
  not KeyNOTGate_0_87(N807, KeyNOTWire_0[87]);
  and AND2_318 (keyinput_Wire_0[199], N219, N802);
  xnor keyGate_0_199(N808, keyinput199, keyinput_Wire_0[199]);
  and AND2_319 (keyinput_Wire_0[200], N219, N803);
  xor keyGate_0_200(N809, keyinput200, keyinput_Wire_0[200]);
  and AND2_320 (keyinput_Wire_0[201], N219, N804);
  xor keyGate_0_201(N810, keyinput201, keyinput_Wire_0[201]);
  nand NAND4_321 (keyinput_Wire_0[202], N805, N787, N731, N529);
  xnor keyGate_0_202(N811, keyinput202, keyinput_Wire_0[202]);
  nand NAND2_322 (keyinput_Wire_0[203], N619, N796);
  xnor keyGate_0_203(N812, keyinput203, keyinput_Wire_0[203]);
  nand NAND3_323 (keyinput_Wire_0[204], N609, N619, N796);
  xor keyGate_0_204(KeyNOTWire_0[88], keyinput204, keyinput_Wire_0[204]);
  not KeyNOTGate_0_88(N813, KeyNOTWire_0[88]);
  nand NAND4_324 (keyinput_Wire_0[205], N600, N609, N619, N796);
  xor keyGate_0_205(N814, keyinput205, keyinput_Wire_0[205]);
  nand NAND4_325 (keyinput_Wire_0[206], N738, N765, N766, N814);
  xor keyGate_0_206(KeyNOTWire_0[89], keyinput206, keyinput_Wire_0[206]);
  not KeyNOTGate_0_89(N815, KeyNOTWire_0[89]);
  nand NAND3_326 (keyinput_Wire_0[207], N741, N764, N813);
  xor keyGate_0_207(N819, keyinput207, keyinput_Wire_0[207]);
  nand NAND2_327 (keyinput_Wire_0[208], N744, N812);
  xor keyGate_0_208(N822, keyinput208, keyinput_Wire_0[208]);
  nor NOR2_328 (keyinput_Wire_0[209], N806, N807);
  xnor keyGate_0_209(KeyNOTWire_0[90], keyinput209, keyinput_Wire_0[209]);
  not KeyNOTGate_0_90(N825, KeyNOTWire_0[90]);
  nor NOR2_329 (keyinput_Wire_0[210], N335, N808);
  xnor keyGate_0_210(N826, keyinput210, keyinput_Wire_0[210]);
  nor NOR2_330 (keyinput_Wire_0[211], N336, N809);
  xor keyGate_0_211(N827, keyinput211, keyinput_Wire_0[211]);
  nor NOR2_331 (keyinput_Wire_0[212], N338, N810);
  xnor keyGate_0_212(KeyNOTWire_0[91], keyinput212, keyinput_Wire_0[212]);
  not KeyNOTGate_0_91(N828, KeyNOTWire_0[91]);
  not NOT1_332 (keyinput_Wire_0[213], N811);
  xnor keyGate_0_213(KeyNOTWire_0[92], keyinput213, keyinput_Wire_0[213]);
  not KeyNOTGate_0_92(N829, KeyNOTWire_0[92]);
  nor NOR2_333 (keyinput_Wire_0[214], N665, N815);
  xnor keyGate_0_214(N830, keyinput214, keyinput_Wire_0[214]);
  and AND2_334 (keyinput_Wire_0[215], N665, N815);
  xor keyGate_0_215(KeyNOTWire_0[93], keyinput215, keyinput_Wire_0[215]);
  not KeyNOTGate_0_93(N831, KeyNOTWire_0[93]);
  nor NOR2_335 (keyinput_Wire_0[216], N673, N819);
  xnor keyGate_0_216(KeyNOTWire_0[94], keyinput216, keyinput_Wire_0[216]);
  not KeyNOTGate_0_94(N832, KeyNOTWire_0[94]);
  and AND2_336 (keyinput_Wire_0[217], N673, N819);
  xor keyGate_0_217(N833, keyinput217, keyinput_Wire_0[217]);
  nor NOR2_337 (keyinput_Wire_0[218], N682, N822);
  xnor keyGate_0_218(KeyNOTWire_0[95], keyinput218, keyinput_Wire_0[218]);
  not KeyNOTGate_0_95(N834, KeyNOTWire_0[95]);
  and AND2_338 (keyinput_Wire_0[219], N682, N822);
  xor keyGate_0_219(KeyNOTWire_0[96], keyinput219, keyinput_Wire_0[219]);
  not KeyNOTGate_0_96(N835, KeyNOTWire_0[96]);
  and AND2_339 (keyinput_Wire_0[220], N219, N825);
  xor keyGate_0_220(N836, keyinput220, keyinput_Wire_0[220]);
  nand NAND3_340 (keyinput_Wire_0[221], N826, N777, N704);
  xnor keyGate_0_221(KeyNOTWire_0[97], keyinput221, keyinput_Wire_0[221]);
  not KeyNOTGate_0_97(N837, KeyNOTWire_0[97]);
  nand NAND4_341 (keyinput_Wire_0[222], N827, N781, N712, N527);
  xnor keyGate_0_222(N838, keyinput222, keyinput_Wire_0[222]);
  nand NAND4_342 (keyinput_Wire_0[223], N828, N785, N721, N528);
  xnor keyGate_0_223(N839, keyinput223, keyinput_Wire_0[223]);
  not NOT1_343 (keyinput_Wire_0[224], N829);
  xor keyGate_0_224(N840, keyinput224, keyinput_Wire_0[224]);
  nand NAND2_344 (keyinput_Wire_0[225], N815, N593);
  xnor keyGate_0_225(KeyNOTWire_0[98], keyinput225, keyinput_Wire_0[225]);
  not KeyNOTGate_0_98(N841, KeyNOTWire_0[98]);
  nor NOR2_345 (keyinput_Wire_0[226], N830, N831);
  xor keyGate_0_226(N842, keyinput226, keyinput_Wire_0[226]);
  nor NOR2_346 (keyinput_Wire_0[227], N832, N833);
  xor keyGate_0_227(N843, keyinput227, keyinput_Wire_0[227]);
  nor NOR2_347 (keyinput_Wire_0[228], N834, N835);
  xnor keyGate_0_228(N844, keyinput228, keyinput_Wire_0[228]);
  nor NOR2_348 (keyinput_Wire_0[229], N334, N836);
  xor keyGate_0_229(KeyNOTWire_0[99], keyinput229, keyinput_Wire_0[229]);
  not KeyNOTGate_0_99(N845, KeyNOTWire_0[99]);
  not NOT1_349 (keyinput_Wire_0[230], N837);
  xor keyGate_0_230(KeyNOTWire_0[100], keyinput230, keyinput_Wire_0[230]);
  not KeyNOTGate_0_100(N846, KeyNOTWire_0[100]);
  not NOT1_350 (keyinput_Wire_0[231], N838);
  xnor keyGate_0_231(KeyNOTWire_0[101], keyinput231, keyinput_Wire_0[231]);
  not KeyNOTGate_0_101(N847, KeyNOTWire_0[101]);
  not NOT1_351 (keyinput_Wire_0[232], N839);
  xnor keyGate_0_232(KeyNOTWire_0[102], keyinput232, keyinput_Wire_0[232]);
  not KeyNOTGate_0_102(N848, KeyNOTWire_0[102]);
  and AND2_352 (keyinput_Wire_0[233], N735, N841);
  xor keyGate_0_233(KeyNOTWire_0[103], keyinput233, keyinput_Wire_0[233]);
  not KeyNOTGate_0_103(N849, KeyNOTWire_0[103]);
buf BUFF1_353 (N850, N840);
  and AND2_354 (keyinput_Wire_0[234], N219, N842);
  xnor keyGate_0_234(N851, keyinput234, keyinput_Wire_0[234]);
  and AND2_355 (keyinput_Wire_0[235], N219, N843);
  xor keyGate_0_235(N852, keyinput235, keyinput_Wire_0[235]);
  and AND2_356 (keyinput_Wire_0[236], N219, N844);
  xnor keyGate_0_236(KeyNOTWire_0[104], keyinput236, keyinput_Wire_0[236]);
  not KeyNOTGate_0_104(N853, KeyNOTWire_0[104]);
  nand NAND3_357 (keyinput_Wire_0[237], N845, N772, N696);
  xor keyGate_0_237(N854, keyinput237, keyinput_Wire_0[237]);
  not NOT1_358 (keyinput_Wire_0[238], N846);
  xor keyGate_0_238(KeyNOTWire_0[105], keyinput238, keyinput_Wire_0[238]);
  not KeyNOTGate_0_105(N855, KeyNOTWire_0[105]);
  not NOT1_359 (keyinput_Wire_0[239], N847);
  xor keyGate_0_239(KeyNOTWire_0[106], keyinput239, keyinput_Wire_0[239]);
  not KeyNOTGate_0_106(N856, KeyNOTWire_0[106]);
  not NOT1_360 (keyinput_Wire_0[240], N848);
  xor keyGate_0_240(N857, keyinput240, keyinput_Wire_0[240]);
  not NOT1_361 (keyinput_Wire_0[241], N849);
  xor keyGate_0_241(KeyNOTWire_0[107], keyinput241, keyinput_Wire_0[241]);
  not KeyNOTGate_0_107(N858, KeyNOTWire_0[107]);
  nor NOR2_362 (keyinput_Wire_0[242], N417, N851);
  xnor keyGate_0_242(N859, keyinput242, keyinput_Wire_0[242]);
  nor NOR2_363 (keyinput_Wire_0[243], N332, N852);
  xor keyGate_0_243(N860, keyinput243, keyinput_Wire_0[243]);
  nor NOR2_364 (keyinput_Wire_0[244], N333, N853);
  xor keyGate_0_244(N861, keyinput244, keyinput_Wire_0[244]);
  not NOT1_365 (keyinput_Wire_0[245], N854);
  xnor keyGate_0_245(KeyNOTWire_0[108], keyinput245, keyinput_Wire_0[245]);
  not KeyNOTGate_0_108(N862, KeyNOTWire_0[108]);
buf BUFF1_366 (N863, N855);
  buf BUFF1_367 (keyinput_Wire_1, N856);
  xor keyGate_1_7(N864, KeyWire_0_2, keyinput_Wire_1);
buf BUFF1_368 (N865, N857);
buf BUFF1_369 (N866, N858);
  nand NAND3_370 (keyinput_Wire_0[246], N859, N769, N669);
  xnor keyGate_0_246(N867, keyinput246, keyinput_Wire_0[246]);
  nand NAND3_371 (keyinput_Wire_0[247], N860, N770, N677);
  xnor keyGate_0_247(N868, keyinput247, keyinput_Wire_0[247]);
  nand NAND3_372 (keyinput_Wire_0[248], N861, N771, N686);
  xor keyGate_0_248(KeyNOTWire_0[109], keyinput248, keyinput_Wire_0[248]);
  not KeyNOTGate_0_109(N869, KeyNOTWire_0[109]);
  not NOT1_373 (keyinput_Wire_0[249], N862);
  xor keyGate_0_249(N870, keyinput249, keyinput_Wire_0[249]);
  not NOT1_374 (keyinput_Wire_0[250], N867);
  xor keyGate_0_250(KeyNOTWire_0[110], keyinput250, keyinput_Wire_0[250]);
  not KeyNOTGate_0_110(N871, KeyNOTWire_0[110]);
  not NOT1_375 (keyinput_Wire_0[251], N868);
  xnor keyGate_0_251(N872, keyinput251, keyinput_Wire_0[251]);
  not NOT1_376 (keyinput_Wire_0[252], N869);
  xnor keyGate_0_252(KeyNOTWire_0[111], keyinput252, keyinput_Wire_0[252]);
  not KeyNOTGate_0_111(N873, KeyNOTWire_0[111]);
buf BUFF1_377 (N874, N870);
  not NOT1_378 (keyinput_Wire_0[253], N871);
  xnor keyGate_0_253(KeyNOTWire_0[112], keyinput253, keyinput_Wire_0[253]);
  not KeyNOTGate_0_112(N875, KeyNOTWire_0[112]);
  not NOT1_379 (keyinput_Wire_0[254], N872);
  xnor keyGate_0_254(N876, keyinput254, keyinput_Wire_0[254]);
  not NOT1_380 (keyinput_Wire_0[255], N873);
  xor keyGate_0_255(KeyNOTWire_0[113], keyinput255, keyinput_Wire_0[255]);
  not KeyNOTGate_0_113(N877, KeyNOTWire_0[113]);
buf BUFF1_381 (N878, N875);
buf BUFF1_382 (N879, N876);
buf BUFF1_383 (N880, N877);

AntiSAT some_name( KeyWire_0_2, N246, N8, N267, N171, N156, N121, N106, N51, N261, N228, N201, N143, N26, N72, N130, N138, N219, N237, N29, N165, N1, N13, N153, N85, N87, N159, N195, N146, N73, N189, N101, N96, N210, N55, N89, N260, N59, N207, N17, N88, N75, N126, N177, N149, N90, N74, N116, N255, N91, N268, N259, N111, N68, N42, N183, N80, N152, N135, N86, N36, keyinput256, keyinput257, keyinput258, keyinput259, keyinput260, keyinput261, keyinput262, keyinput263, keyinput264, keyinput265, keyinput266, keyinput267, keyinput268, keyinput269, keyinput270, keyinput271, keyinput272, keyinput273, keyinput274, keyinput275, keyinput276, keyinput277, keyinput278, keyinput279, keyinput280, keyinput281, keyinput282, keyinput283, keyinput284, keyinput285, keyinput286, keyinput287, keyinput288, keyinput289, keyinput290, keyinput291, keyinput292, keyinput293, keyinput294, keyinput295, keyinput296, keyinput297, keyinput298, keyinput299, keyinput300, keyinput301, keyinput302, keyinput303, keyinput304, keyinput305, keyinput306, keyinput307, keyinput308, keyinput309, keyinput310, keyinput311, keyinput312, keyinput313, keyinput314, keyinput315, keyinput316, keyinput317, keyinput318, keyinput319, keyinput320, keyinput321, keyinput322, keyinput323, keyinput324, keyinput325, keyinput326, keyinput327, keyinput328, keyinput329, keyinput330, keyinput331, keyinput332, keyinput333, keyinput334, keyinput335, keyinput336, keyinput337, keyinput338, keyinput339, keyinput340, keyinput341, keyinput342, keyinput343, keyinput344, keyinput345, keyinput346, keyinput347, keyinput348, keyinput349, keyinput350, keyinput351, keyinput352, keyinput353, keyinput354, keyinput355, keyinput356, keyinput357, keyinput358, keyinput359, keyinput360, keyinput361, keyinput362, keyinput363, keyinput364, keyinput365, keyinput366, keyinput367, keyinput368, keyinput369, keyinput370, keyinput371, keyinput372, keyinput373, keyinput374, keyinput375,
       keyinput376, keyinput377, keyinput378, keyinput379, keyinput380,
       keyinput381, keyinput382, keyinput383, keyinput384, keyinput385,
       keyinput386, keyinput387, keyinput388, keyinput389, keyinput390,
       keyinput391, keyinput392, keyinput393, keyinput394, keyinput395,
       keyinput396, keyinput397, keyinput398, keyinput399, keyinput400,
       keyinput401, keyinput402, keyinput403, keyinput404, keyinput405,
       keyinput406, keyinput407, keyinput408, keyinput409, keyinput410,
       keyinput411, keyinput412, keyinput413, keyinput414, keyinput415,
       keyinput416, keyinput417, keyinput418, keyinput419, keyinput420,
       keyinput421, keyinput422, keyinput423, keyinput424, keyinput425,
       keyinput426, keyinput427, keyinput428, keyinput429, keyinput430,
       keyinput431, keyinput432, keyinput433, keyinput434, keyinput435);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N246, N8, N267, N171, N156, N121, N106, N51, N261, N228, N201, N143, N26, N72, N130, N138, N219, N237, N29, N165, N1, N13, N153, N85, N87, N159, N195, N146, N73, N189, N101, N96, N210, N55, N89, N260, N59, N207, N17, N88, N75, N126, N177, N149, N90, N74, N116, N255, N91, N268, N259, N111, N68, N42, N183, N80, N152, N135, N86, N36, keyinput256, keyinput257, keyinput258, keyinput259, keyinput260, keyinput261, keyinput262, keyinput263, keyinput264, keyinput265, keyinput266, keyinput267, keyinput268, keyinput269, keyinput270, keyinput271, keyinput272, keyinput273, keyinput274, keyinput275, keyinput276, keyinput277, keyinput278, keyinput279, keyinput280, keyinput281, keyinput282, keyinput283, keyinput284, keyinput285, keyinput286, keyinput287, keyinput288, keyinput289, keyinput290, keyinput291, keyinput292, keyinput293, keyinput294, keyinput295, keyinput296, keyinput297, keyinput298, keyinput299, keyinput300, keyinput301, keyinput302, keyinput303, keyinput304, keyinput305, keyinput306, keyinput307, keyinput308, keyinput309, keyinput310, keyinput311, keyinput312, keyinput313, keyinput314, keyinput315, keyinput316, keyinput317, keyinput318, keyinput319, keyinput320, keyinput321, keyinput322, keyinput323, keyinput324, keyinput325, keyinput326, keyinput327, keyinput328, keyinput329, keyinput330, keyinput331, keyinput332, keyinput333, keyinput334, keyinput335, keyinput336, keyinput337, keyinput338, keyinput339, keyinput340, keyinput341, keyinput342, keyinput343, keyinput344, keyinput345, keyinput346, keyinput347, keyinput348, keyinput349, keyinput350, keyinput351, keyinput352, keyinput353, keyinput354, keyinput355, keyinput356, keyinput357, keyinput358, keyinput359, keyinput360, keyinput361, keyinput362, keyinput363, keyinput364, keyinput365, keyinput366, keyinput367, keyinput368, keyinput369, keyinput370, keyinput371, keyinput372, keyinput373, keyinput374, keyinput375 ,
        keyinput376, keyinput377, keyinput378, keyinput379, keyinput380,
        keyinput381, keyinput382, keyinput383, keyinput384, keyinput385,
        keyinput386, keyinput387, keyinput388, keyinput389, keyinput390,
        keyinput391, keyinput392, keyinput393, keyinput394, keyinput395,
        keyinput396, keyinput397, keyinput398, keyinput399, keyinput400,
        keyinput401, keyinput402, keyinput403, keyinput404, keyinput405,
        keyinput406, keyinput407, keyinput408, keyinput409, keyinput410,
        keyinput411, keyinput412, keyinput413, keyinput414, keyinput415,
        keyinput416, keyinput417, keyinput418, keyinput419, keyinput420,
        keyinput421, keyinput422, keyinput423, keyinput424, keyinput425,
        keyinput426, keyinput427, keyinput428, keyinput429, keyinput430,
        keyinput431, keyinput432, keyinput433, keyinput434, keyinput435);

  input keyinput376, keyinput377, keyinput378, keyinput379, keyinput380;
  input keyinput381, keyinput382, keyinput383, keyinput384, keyinput385;
  input keyinput386, keyinput387, keyinput388, keyinput389, keyinput390;
  input keyinput391, keyinput392, keyinput393, keyinput394, keyinput395;
  input keyinput396, keyinput397, keyinput398, keyinput399, keyinput400;
  input keyinput401, keyinput402, keyinput403, keyinput404, keyinput405;
  input keyinput406, keyinput407, keyinput408, keyinput409, keyinput410;
  input keyinput411, keyinput412, keyinput413, keyinput414, keyinput415;
  input keyinput416, keyinput417, keyinput418, keyinput419, keyinput420;
  input keyinput421, keyinput422, keyinput423, keyinput424, keyinput425;
  input keyinput426, keyinput427, keyinput428, keyinput429, keyinput430;
  input keyinput431, keyinput432, keyinput433, keyinput434, keyinput435;

  wire [0:59] keyNTin_Wire_1;
  wire [0:26] KeyNOTWire_1;

  input N246, N8, N267, N171, N156, N121, N106, N51, N261, N228, N201, N143, N26, N72, N130, N138, N219, N237, N29, N165, N1, N13, N153, N85, N87, N159, N195, N146, N73, N189, N101, N96, N210, N55, N89, N260, N59, N207, N17, N88, N75, N126, N177, N149, N90, N74, N116, N255, N91, N268, N259, N111, N68, N42, N183, N80, N152, N135, N86, N36;
  input keyinput256, keyinput257, keyinput258, keyinput259, keyinput260, keyinput261, keyinput262, keyinput263, keyinput264, keyinput265, keyinput266, keyinput267, keyinput268, keyinput269, keyinput270, keyinput271, keyinput272, keyinput273, keyinput274, keyinput275, keyinput276, keyinput277, keyinput278, keyinput279, keyinput280, keyinput281, keyinput282, keyinput283, keyinput284, keyinput285, keyinput286, keyinput287, keyinput288, keyinput289, keyinput290, keyinput291, keyinput292, keyinput293, keyinput294, keyinput295, keyinput296, keyinput297, keyinput298, keyinput299, keyinput300, keyinput301, keyinput302, keyinput303, keyinput304, keyinput305, keyinput306, keyinput307, keyinput308, keyinput309, keyinput310, keyinput311, keyinput312, keyinput313, keyinput314, keyinput315, keyinput316, keyinput317, keyinput318, keyinput319, keyinput320, keyinput321, keyinput322, keyinput323, keyinput324, keyinput325, keyinput326, keyinput327, keyinput328, keyinput329, keyinput330, keyinput331, keyinput332, keyinput333, keyinput334, keyinput335, keyinput336, keyinput337, keyinput338, keyinput339, keyinput340, keyinput341, keyinput342, keyinput343, keyinput344, keyinput345, keyinput346, keyinput347, keyinput348, keyinput349, keyinput350, keyinput351, keyinput352, keyinput353, keyinput354, keyinput355, keyinput356, keyinput357, keyinput358, keyinput359, keyinput360, keyinput361, keyinput362, keyinput363, keyinput364, keyinput365, keyinput366, keyinput367, keyinput368, keyinput369, keyinput370, keyinput371, keyinput372, keyinput373, keyinput374, keyinput375;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83, newWire_84, newWire_85, newWire_86, newWire_87, newWire_88, newWire_89, newWire_90, newWire_91, newWire_92, newWire_93, newWire_94, newWire_95, newWire_96, newWire_97, newWire_98, newWire_99, newWire_100, newWire_101, newWire_102, newWire_103, newWire_104, newWire_105, newWire_106, newWire_107, newWire_108, newWire_109, newWire_110, newWire_111, newWire_112, newWire_113, newWire_114, newWire_115, newWire_116, newWire_117, newWire_118, newWire_119, newWire_120, newWire_121 ;

  xnor KeyGate0 (keyNTin_Wire_1[0], N246, keyinput256);
  xnor keyNTinGate_1_0(newWire_0, keyinput376, keyNTin_Wire_1[0]);
  xor  KeyGate1 (newWire_1, N8, keyinput257);
  xor  KeyGate2 (newWire_2, N267, keyinput258);
  xor  KeyGate3 (keyNTin_Wire_1[1], N171, keyinput259);
  xnor keyNTinGate_1_1(newWire_3, keyinput377, keyNTin_Wire_1[1]);
  xnor KeyGate4 (keyNTin_Wire_1[2], N156, keyinput260);
  xnor keyNTinGate_1_2(KeyNOTWire_1[0], keyinput378, keyNTin_Wire_1[2]);
  not KeyNOTGate_1_0(newWire_4, KeyNOTWire_1[0]);
  xor  KeyGate5 (keyNTin_Wire_1[3], N121, keyinput261);
  xnor keyNTinGate_1_3(newWire_5, keyinput379, keyNTin_Wire_1[3]);
  xor  KeyGate6 (newWire_6, N106, keyinput262);
  xor  KeyGate7 (keyNTin_Wire_1[4], N51, keyinput263);
  xor keyNTinGate_1_4(newWire_7, keyinput380, keyNTin_Wire_1[4]);
  xnor KeyGate8 (keyNTin_Wire_1[5], N261, keyinput264);
  xnor keyNTinGate_1_5(newWire_8, keyinput381, keyNTin_Wire_1[5]);
  xor  KeyGate9 (keyNTin_Wire_1[6], N228, keyinput265);
  xnor keyNTinGate_1_6(KeyNOTWire_1[1], keyinput382, keyNTin_Wire_1[6]);
  not KeyNOTGate_1_1(newWire_9, KeyNOTWire_1[1]);
  xor  KeyGate10 (newWire_10, N201, keyinput266);
  xnor KeyGate11 (newWire_11, N143, keyinput267);
  xnor KeyGate12 (keyNTin_Wire_1[7], N26, keyinput268);
  xnor keyNTinGate_1_7(KeyNOTWire_1[2], keyinput383, keyNTin_Wire_1[7]);
  not KeyNOTGate_1_2(newWire_12, KeyNOTWire_1[2]);
  xnor KeyGate13 (newWire_13, N72, keyinput269);
  xnor KeyGate14 (newWire_14, N130, keyinput270);
  xor  KeyGate15 (keyNTin_Wire_1[8], N138, keyinput271);
  xor keyNTinGate_1_8(KeyNOTWire_1[3], keyinput384, keyNTin_Wire_1[8]);
  not KeyNOTGate_1_3(newWire_15, KeyNOTWire_1[3]);
  xnor KeyGate16 (keyNTin_Wire_1[9], N219, keyinput272);
  xnor keyNTinGate_1_9(KeyNOTWire_1[4], keyinput385, keyNTin_Wire_1[9]);
  not KeyNOTGate_1_4(newWire_16, KeyNOTWire_1[4]);
  xnor KeyGate17 (newWire_17, N237, keyinput273);
  xor  KeyGate18 (keyNTin_Wire_1[10], N29, keyinput274);
  xor keyNTinGate_1_10(KeyNOTWire_1[5], keyinput386, keyNTin_Wire_1[10]);
  not KeyNOTGate_1_5(newWire_18, KeyNOTWire_1[5]);
  xor  KeyGate19 (newWire_19, N165, keyinput275);
  xor  KeyGate20 (keyNTin_Wire_1[11], N1, keyinput276);
  xor keyNTinGate_1_11(KeyNOTWire_1[6], keyinput387, keyNTin_Wire_1[11]);
  not KeyNOTGate_1_6(newWire_20, KeyNOTWire_1[6]);
  xor  KeyGate21 (newWire_21, N13, keyinput277);
  xnor KeyGate22 (newWire_22, N153, keyinput278);
  xnor KeyGate23 (keyNTin_Wire_1[12], N85, keyinput279);
  xnor keyNTinGate_1_12(KeyNOTWire_1[7], keyinput388, keyNTin_Wire_1[12]);
  not KeyNOTGate_1_7(newWire_23, KeyNOTWire_1[7]);
  xnor KeyGate24 (keyNTin_Wire_1[13], N87, keyinput280);
  xor keyNTinGate_1_13(newWire_24, keyinput389, keyNTin_Wire_1[13]);
  xor  KeyGate25 (newWire_25, N159, keyinput281);
  xnor KeyGate26 (keyNTin_Wire_1[14], N195, keyinput282);
  xnor keyNTinGate_1_14(newWire_26, keyinput390, keyNTin_Wire_1[14]);
  xnor KeyGate27 (newWire_27, N146, keyinput283);
  xor  KeyGate28 (keyNTin_Wire_1[15], N73, keyinput284);
  xnor keyNTinGate_1_15(KeyNOTWire_1[8], keyinput391, keyNTin_Wire_1[15]);
  not KeyNOTGate_1_8(newWire_28, KeyNOTWire_1[8]);
  xor  KeyGate29 (keyNTin_Wire_1[16], N189, keyinput285);
  xnor keyNTinGate_1_16(newWire_29, keyinput392, keyNTin_Wire_1[16]);
  xor  KeyGate30 (newWire_30, N101, keyinput286);
  xor  KeyGate31 (newWire_31, N96, keyinput287);
  xnor KeyGate32 (keyNTin_Wire_1[17], N210, keyinput288);
  xor keyNTinGate_1_17(KeyNOTWire_1[9], keyinput393, keyNTin_Wire_1[17]);
  not KeyNOTGate_1_9(newWire_32, KeyNOTWire_1[9]);
  xnor KeyGate33 (newWire_33, N55, keyinput289);
  xor  KeyGate34 (newWire_34, N89, keyinput290);
  xnor KeyGate35 (newWire_35, N260, keyinput291);
  xor  KeyGate36 (newWire_36, N59, keyinput292);
  xor  KeyGate37 (newWire_37, N207, keyinput293);
  xnor KeyGate38 (newWire_38, N17, keyinput294);
  xor  KeyGate39 (newWire_39, N88, keyinput295);
  xnor KeyGate40 (keyNTin_Wire_1[18], N75, keyinput296);
  xnor keyNTinGate_1_18(newWire_40, keyinput394, keyNTin_Wire_1[18]);
  xor  KeyGate41 (newWire_41, N126, keyinput297);
  xor  KeyGate42 (keyNTin_Wire_1[19], N177, keyinput298);
  xor keyNTinGate_1_19(KeyNOTWire_1[10], keyinput395, keyNTin_Wire_1[19]);
  not KeyNOTGate_1_10(newWire_42, KeyNOTWire_1[10]);
  xnor KeyGate43 (keyNTin_Wire_1[20], N149, keyinput299);
  xnor keyNTinGate_1_20(KeyNOTWire_1[11], keyinput396, keyNTin_Wire_1[20]);
  not KeyNOTGate_1_11(newWire_43, KeyNOTWire_1[11]);
  xor  KeyGate44 (newWire_44, N90, keyinput300);
  xor  KeyGate45 (newWire_45, N74, keyinput301);
  xnor KeyGate46 (newWire_46, N116, keyinput302);
  xor  KeyGate47 (newWire_47, N255, keyinput303);
  xor  KeyGate48 (keyNTin_Wire_1[21], N91, keyinput304);
  xnor keyNTinGate_1_21(KeyNOTWire_1[12], keyinput397, keyNTin_Wire_1[21]);
  not KeyNOTGate_1_12(newWire_48, KeyNOTWire_1[12]);
  xor  KeyGate49 (keyNTin_Wire_1[22], N268, keyinput305);
  xor keyNTinGate_1_22(newWire_49, keyinput398, keyNTin_Wire_1[22]);
  xor  KeyGate50 (keyNTin_Wire_1[23], N259, keyinput306);
  xor keyNTinGate_1_23(newWire_50, keyinput399, keyNTin_Wire_1[23]);
  xnor KeyGate51 (newWire_51, N111, keyinput307);
  xnor KeyGate52 (keyNTin_Wire_1[24], N68, keyinput308);
  xor keyNTinGate_1_24(newWire_52, keyinput400, keyNTin_Wire_1[24]);
  xnor KeyGate53 (keyNTin_Wire_1[25], N42, keyinput309);
  xnor keyNTinGate_1_25(KeyNOTWire_1[13], keyinput401, keyNTin_Wire_1[25]);
  not KeyNOTGate_1_13(newWire_53, KeyNOTWire_1[13]);
  xor  KeyGate54 (keyNTin_Wire_1[26], N183, keyinput310);
  xnor keyNTinGate_1_26(KeyNOTWire_1[14], keyinput402, keyNTin_Wire_1[26]);
  not KeyNOTGate_1_14(newWire_54, KeyNOTWire_1[14]);
  xor  KeyGate55 (keyNTin_Wire_1[27], N80, keyinput311);
  xor keyNTinGate_1_27(newWire_55, keyinput403, keyNTin_Wire_1[27]);
  xor  KeyGate56 (newWire_56, N152, keyinput312);
  xnor KeyGate57 (newWire_57, N135, keyinput313);
  xor  KeyGate58 (keyNTin_Wire_1[28], N86, keyinput314);
  xnor keyNTinGate_1_28(KeyNOTWire_1[15], keyinput404, keyNTin_Wire_1[28]);
  not KeyNOTGate_1_15(newWire_58, KeyNOTWire_1[15]);
  xnor KeyGate59 (newWire_59, N36, keyinput315);
  xnor KeyGate60 (newWire_60, N246, keyinput316);
  xnor KeyGate61 (newWire_61, N8, keyinput317);
  xor  KeyGate62 (newWire_62, N267, keyinput318);
  xnor KeyGate63 (newWire_63, N171, keyinput319);
  xor  KeyGate64 (keyNTin_Wire_1[29], N156, keyinput320);
  xor keyNTinGate_1_29(KeyNOTWire_1[16], keyinput405, keyNTin_Wire_1[29]);
  not KeyNOTGate_1_16(newWire_64, KeyNOTWire_1[16]);
  xor  KeyGate65 (newWire_65, N121, keyinput321);
  xnor KeyGate66 (newWire_66, N106, keyinput322);
  xnor KeyGate67 (keyNTin_Wire_1[30], N51, keyinput323);
  xor keyNTinGate_1_30(KeyNOTWire_1[17], keyinput406, keyNTin_Wire_1[30]);
  not KeyNOTGate_1_17(newWire_67, KeyNOTWire_1[17]);
  xnor KeyGate68 (keyNTin_Wire_1[31], N261, keyinput324);
  xnor keyNTinGate_1_31(newWire_68, keyinput407, keyNTin_Wire_1[31]);
  xor  KeyGate69 (keyNTin_Wire_1[32], N228, keyinput325);
  xnor keyNTinGate_1_32(KeyNOTWire_1[18], keyinput408, keyNTin_Wire_1[32]);
  not KeyNOTGate_1_18(newWire_69, KeyNOTWire_1[18]);
  xor  KeyGate70 (keyNTin_Wire_1[33], N201, keyinput326);
  xor keyNTinGate_1_33(KeyNOTWire_1[19], keyinput409, keyNTin_Wire_1[33]);
  not KeyNOTGate_1_19(newWire_70, KeyNOTWire_1[19]);
  xnor KeyGate71 (keyNTin_Wire_1[34], N143, keyinput327);
  xor keyNTinGate_1_34(KeyNOTWire_1[20], keyinput410, keyNTin_Wire_1[34]);
  not KeyNOTGate_1_20(newWire_71, KeyNOTWire_1[20]);
  xor  KeyGate72 (keyNTin_Wire_1[35], N26, keyinput328);
  xnor keyNTinGate_1_35(newWire_72, keyinput411, keyNTin_Wire_1[35]);
  xnor KeyGate73 (newWire_73, N72, keyinput329);
  xor  KeyGate74 (keyNTin_Wire_1[36], N130, keyinput330);
  xnor keyNTinGate_1_36(newWire_74, keyinput412, keyNTin_Wire_1[36]);
  xor  KeyGate75 (newWire_75, N138, keyinput331);
  xnor KeyGate76 (newWire_76, N219, keyinput332);
  xnor KeyGate77 (newWire_77, N237, keyinput333);
  xnor KeyGate78 (newWire_78, N29, keyinput334);
  xor  KeyGate79 (newWire_79, N165, keyinput335);
  xnor KeyGate80 (keyNTin_Wire_1[37], N1, keyinput336);
  xor keyNTinGate_1_37(newWire_80, keyinput413, keyNTin_Wire_1[37]);
  xnor KeyGate81 (newWire_81, N13, keyinput337);
  xnor KeyGate82 (newWire_82, N153, keyinput338);
  xnor KeyGate83 (keyNTin_Wire_1[38], N85, keyinput339);
  xor keyNTinGate_1_38(KeyNOTWire_1[21], keyinput414, keyNTin_Wire_1[38]);
  not KeyNOTGate_1_21(newWire_83, KeyNOTWire_1[21]);
  xor  KeyGate84 (keyNTin_Wire_1[39], N87, keyinput340);
  xnor keyNTinGate_1_39(KeyNOTWire_1[22], keyinput415, keyNTin_Wire_1[39]);
  not KeyNOTGate_1_22(newWire_84, KeyNOTWire_1[22]);
  xnor KeyGate85 (newWire_85, N159, keyinput341);
  xnor KeyGate86 (newWire_86, N195, keyinput342);
  xnor KeyGate87 (keyNTin_Wire_1[40], N146, keyinput343);
  xor keyNTinGate_1_40(newWire_87, keyinput416, keyNTin_Wire_1[40]);
  xor  KeyGate88 (keyNTin_Wire_1[41], N73, keyinput344);
  xnor keyNTinGate_1_41(KeyNOTWire_1[23], keyinput417, keyNTin_Wire_1[41]);
  not KeyNOTGate_1_23(newWire_88, KeyNOTWire_1[23]);
  xnor KeyGate89 (newWire_89, N189, keyinput345);
  xor  KeyGate90 (keyNTin_Wire_1[42], N101, keyinput346);
  xnor keyNTinGate_1_42(newWire_90, keyinput418, keyNTin_Wire_1[42]);
  xor  KeyGate91 (keyNTin_Wire_1[43], N96, keyinput347);
  xnor keyNTinGate_1_43(KeyNOTWire_1[24], keyinput419, keyNTin_Wire_1[43]);
  not KeyNOTGate_1_24(newWire_91, KeyNOTWire_1[24]);
  xor  KeyGate92 (keyNTin_Wire_1[44], N210, keyinput348);
  xor keyNTinGate_1_44(newWire_92, keyinput420, keyNTin_Wire_1[44]);
  xnor KeyGate93 (newWire_93, N55, keyinput349);
  xor  KeyGate94 (newWire_94, N89, keyinput350);
  xor  KeyGate95 (keyNTin_Wire_1[45], N260, keyinput351);
  xnor keyNTinGate_1_45(newWire_95, keyinput421, keyNTin_Wire_1[45]);
  xnor KeyGate96 (keyNTin_Wire_1[46], N59, keyinput352);
  xor keyNTinGate_1_46(newWire_96, keyinput422, keyNTin_Wire_1[46]);
  xor  KeyGate97 (keyNTin_Wire_1[47], N207, keyinput353);
  xnor keyNTinGate_1_47(newWire_97, keyinput423, keyNTin_Wire_1[47]);
  xnor KeyGate98 (keyNTin_Wire_1[48], N17, keyinput354);
  xnor keyNTinGate_1_48(newWire_98, keyinput424, keyNTin_Wire_1[48]);
  xnor KeyGate99 (newWire_99, N88, keyinput355);
  xnor KeyGate100 (newWire_100, N75, keyinput356);
  xnor KeyGate101 (newWire_101, N126, keyinput357);
  xnor KeyGate102 (newWire_102, N177, keyinput358);
  xnor KeyGate103 (newWire_103, N149, keyinput359);
  xor  KeyGate104 (keyNTin_Wire_1[49], N90, keyinput360);
  xnor keyNTinGate_1_49(KeyNOTWire_1[25], keyinput425, keyNTin_Wire_1[49]);
  not KeyNOTGate_1_25(newWire_104, KeyNOTWire_1[25]);
  xnor KeyGate105 (newWire_105, N74, keyinput361);
  xnor KeyGate106 (newWire_106, N116, keyinput362);
  xnor KeyGate107 (keyNTin_Wire_1[50], N255, keyinput363);
  xnor keyNTinGate_1_50(newWire_107, keyinput426, keyNTin_Wire_1[50]);
  xnor KeyGate108 (keyNTin_Wire_1[51], N91, keyinput364);
  xor keyNTinGate_1_51(newWire_108, keyinput427, keyNTin_Wire_1[51]);
  xnor KeyGate109 (keyNTin_Wire_1[52], N268, keyinput365);
  xor keyNTinGate_1_52(newWire_109, keyinput428, keyNTin_Wire_1[52]);
  xor  KeyGate110 (keyNTin_Wire_1[53], N259, keyinput366);
  xor keyNTinGate_1_53(newWire_110, keyinput429, keyNTin_Wire_1[53]);
  xnor KeyGate111 (keyNTin_Wire_1[54], N111, keyinput367);
  xnor keyNTinGate_1_54(KeyNOTWire_1[26], keyinput430, keyNTin_Wire_1[54]);
  not KeyNOTGate_1_26(newWire_111, KeyNOTWire_1[26]);
  xnor KeyGate112 (newWire_112, N68, keyinput368);
  xor  KeyGate113 (newWire_113, N42, keyinput369);
  xnor KeyGate114 (newWire_114, N183, keyinput370);
  xnor KeyGate115 (newWire_115, N80, keyinput371);
  xor  KeyGate116 (keyNTin_Wire_1[55], N152, keyinput372);
  xnor keyNTinGate_1_55(newWire_116, keyinput431, keyNTin_Wire_1[55]);
  xor  KeyGate117 (keyNTin_Wire_1[56], N135, keyinput373);
  xor keyNTinGate_1_56(newWire_117, keyinput432, keyNTin_Wire_1[56]);
  xor  KeyGate118 (newWire_118, N86, keyinput374);
  xor  KeyGate119 (keyNTin_Wire_1[57], N36, keyinput375);
  xnor keyNTinGate_1_57(newWire_119, keyinput433, keyNTin_Wire_1[57]);
  and some_function (keyNTin_Wire_1[58], newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59 );
  xor keyNTinGate_1_58(newWire_120, keyinput434, keyNTin_Wire_1[58]);
  nand compl_function (keyNTin_Wire_1[59], newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83, newWire_84, newWire_85, newWire_86, newWire_87, newWire_88, newWire_89, newWire_90, newWire_91, newWire_92, newWire_93, newWire_94, newWire_95, newWire_96, newWire_97, newWire_98, newWire_99, newWire_100, newWire_101, newWire_102, newWire_103, newWire_104, newWire_105, newWire_106, newWire_107, newWire_108, newWire_109, newWire_110, newWire_111, newWire_112, newWire_113, newWire_114, newWire_115, newWire_116, newWire_117, newWire_118, newWire_119);
  xor keyNTinGate_1_59(newWire_121, keyinput435, keyNTin_Wire_1[59]);
  and finalAND (KeyWire_0_2, newWire_120, newWire_121);

endmodule /* AntiSAT */
