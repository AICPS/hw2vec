`timescale 1ns / 1ps
// Verilog
// c499
// Ninputs 41
// Noutputs 32
// NtotalGates 202
// XOR2 104
// AND2 40
// NOT1 40
// AND4 8
// OR4 2
// AND5 8

module top (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
                  N753,N754,N755,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
                  keyinput30, keyinput31,
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36,
        keyinput37, keyinput38, keyinput39, keyinput40, keyinput41,
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46,
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51,
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56,
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61,
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66,
        keyinput67, keyinput68, keyinput69, keyinput70, keyinput71,
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76,
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81,
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86,
        keyinput87, keyinput88, keyinput89, keyinput90, keyinput91,
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96,
        keyinput97, keyinput98, keyinput99, keyinput100, keyinput101,
        keyinput102, keyinput103, keyinput104, keyinput105, keyinput106,
        keyinput107, keyinput108, keyinput109, keyinput110, keyinput111,
                  keyinput112, keyinput113,
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
        keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
        keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
        keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
        keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
        keyinput144, keyinput145, keyinput146, keyinput147, keyinput148,
        keyinput149, keyinput150, keyinput151, keyinput152, keyinput153,
        keyinput154);

  input keyinput114, keyinput115, keyinput116, keyinput117, keyinput118;
  input keyinput119, keyinput120, keyinput121, keyinput122, keyinput123;
  input keyinput124, keyinput125, keyinput126, keyinput127, keyinput128;
  input keyinput129, keyinput130, keyinput131, keyinput132, keyinput133;
  input keyinput134, keyinput135, keyinput136, keyinput137, keyinput138;
  input keyinput139, keyinput140, keyinput141, keyinput142, keyinput143;
  input keyinput144, keyinput145, keyinput146, keyinput147, keyinput148;
  input keyinput149, keyinput150, keyinput151, keyinput152, keyinput153;
  input keyinput154;


  input keyinput32, keyinput33, keyinput34, keyinput35, keyinput36;
  input keyinput37, keyinput38, keyinput39, keyinput40, keyinput41;
  input keyinput42, keyinput43, keyinput44, keyinput45, keyinput46;
  input keyinput47, keyinput48, keyinput49, keyinput50, keyinput51;
  input keyinput52, keyinput53, keyinput54, keyinput55, keyinput56;
  input keyinput57, keyinput58, keyinput59, keyinput60, keyinput61;
  input keyinput62, keyinput63, keyinput64, keyinput65, keyinput66;
  input keyinput67, keyinput68, keyinput69, keyinput70, keyinput71;
  input keyinput72, keyinput73, keyinput74, keyinput75, keyinput76;
  input keyinput77, keyinput78, keyinput79, keyinput80, keyinput81;
  input keyinput82, keyinput83, keyinput84, keyinput85, keyinput86;
  input keyinput87, keyinput88, keyinput89, keyinput90, keyinput91;
  input keyinput92, keyinput93, keyinput94, keyinput95, keyinput96;
  input keyinput97, keyinput98, keyinput99, keyinput100, keyinput101;
  input keyinput102, keyinput103, keyinput104, keyinput105, keyinput106;
  input keyinput107, keyinput108, keyinput109, keyinput110, keyinput111;
  input keyinput112, keyinput113;

  wire KeyWire_0_1 , KeyWire_0_2;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31;

  wire [0:31] keyinput_Wire_0;
  wire [0:15] KeyNOTWire_0;

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;

output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723;

xor XOR2_1 (N250, N1, N5);
xor XOR2_2 (N251, N9, N13);
xor XOR2_3 (N252, N17, N21);
xor XOR2_4 (N253, N25, N29);
  xor XOR2_5 (keyinput_Wire_0[0], N33, N37);
  xor keyGate_0_0(N254, keyinput0, keyinput_Wire_0[0]);
xor XOR2_6 (N255, N41, N45);
xor XOR2_7 (N256, N49, N53);
xor XOR2_8 (N257, N57, N61);
xor XOR2_9 (N258, N65, N69);
xor XOR2_10 (N259, N73, N77);
xor XOR2_11 (N260, N81, N85);
xor XOR2_12 (N261, N89, N93);
xor XOR2_13 (N262, N97, N101);
xor XOR2_14 (N263, N105, N109);
xor XOR2_15 (N264, N113, N117);
xor XOR2_16 (N265, N121, N125);
and AND2_17 (N266, N129, N137);
and AND2_18 (N267, N130, N137);
  and AND2_19 (keyinput_Wire_0[1], N131, N137);
  xor keyGate_0_1(KeyNOTWire_0[0], keyinput1, keyinput_Wire_0[1]);
  not KeyNOTGate_0_0(N268, KeyNOTWire_0[0]);
  and AND2_20 (keyinput_Wire_0[2], N132, N137);
  xnor keyGate_0_2(N269, keyinput2, keyinput_Wire_0[2]);
and AND2_21 (N270, N133, N137);
and AND2_22 (N271, N134, N137);
and AND2_23 (N272, N135, N137);
and AND2_24 (N273, N136, N137);
xor XOR2_25 (N274, N1, N17);
  xor XOR2_26 (keyinput_Wire_0[3], N33, N49);
  xor keyGate_0_3(N275, keyinput3, keyinput_Wire_0[3]);
xor XOR2_27 (N276, N5, N21);
xor XOR2_28 (N277, N37, N53);
xor XOR2_29 (N278, N9, N25);
xor XOR2_30 (N279, N41, N57);
xor XOR2_31 (N280, N13, N29);
xor XOR2_32 (N281, N45, N61);
  xor XOR2_33 (keyinput_Wire_0[4], N65, N81);
  xor keyGate_0_4(N282, keyinput4, keyinput_Wire_0[4]);
xor XOR2_34 (N283, N97, N113);
xor XOR2_35 (N284, N69, N85);
xor XOR2_36 (N285, N101, N117);
xor XOR2_37 (N286, N73, N89);
xor XOR2_38 (N287, N105, N121);
xor XOR2_39 (N288, N77, N93);
xor XOR2_40 (N289, N109, N125);
  xor XOR2_41 (keyinput_Wire_0[5], N250, N251);
  xor keyGate_0_5(N290, keyinput5, keyinput_Wire_0[5]);
xor XOR2_42 (N293, N252, N253);
xor XOR2_43 (N296, N254, N255);
  xor XOR2_44 (keyinput_Wire_0[6], N256, N257);
  xor keyGate_0_6(KeyNOTWire_0[1], keyinput6, keyinput_Wire_0[6]);
  not KeyNOTGate_0_1(N299, KeyNOTWire_0[1]);
xor XOR2_45 (N302, N258, N259);
xor XOR2_46 (N305, N260, N261);
xor XOR2_47 (N308, N262, N263);
xor XOR2_48 (N311, N264, N265);
xor XOR2_49 (N314, N274, N275);
  xor XOR2_50 (keyinput_Wire_0[7], N276, N277);
  xnor keyGate_0_7(KeyNOTWire_0[2], keyinput7, keyinput_Wire_0[7]);
  not KeyNOTGate_0_2(N315, KeyNOTWire_0[2]);
xor XOR2_51 (N316, N278, N279);
xor XOR2_52 (N317, N280, N281);
  xor XOR2_53 (keyinput_Wire_0[8], N282, N283);
  xor keyGate_0_8(N318, keyinput8, keyinput_Wire_0[8]);
xor XOR2_54 (N319, N284, N285);
xor XOR2_55 (N320, N286, N287);
xor XOR2_56 (N321, N288, N289);
xor XOR2_57 (N338, N290, N293);
xor XOR2_58 (N339, N296, N299);
xor XOR2_59 (N340, N290, N296);
xor XOR2_60 (N341, N293, N299);
xor XOR2_61 (N342, N302, N305);
xor XOR2_62 (N343, N308, N311);
xor XOR2_63 (N344, N302, N308);
xor XOR2_64 (N345, N305, N311);
xor XOR2_65 (N346, N266, N342);
xor XOR2_66 (N347, N267, N343);
xor XOR2_67 (N348, N268, N344);
  xor XOR2_68 (keyinput_Wire_0[9], N269, N345);
  xor keyGate_0_9(KeyNOTWire_0[3], keyinput9, keyinput_Wire_0[9]);
  not KeyNOTGate_0_3(N349, KeyNOTWire_0[3]);
  xor XOR2_69 (keyinput_Wire_0[10], N270, N338);
  xnor keyGate_0_10(KeyNOTWire_0[4], keyinput10, keyinput_Wire_0[10]);
  not KeyNOTGate_0_4(N350, KeyNOTWire_0[4]);
xor XOR2_70 (N351, N271, N339);
xor XOR2_71 (N352, N272, N340);
  xor XOR2_72 (keyinput_Wire_0[11], N273, N341);
  xor keyGate_0_11(N353, keyinput11, keyinput_Wire_0[11]);
xor XOR2_73 (N354, N314, N346);
xor XOR2_74 (N367, N315, N347);
xor XOR2_75 (N380, N316, N348);
xor XOR2_76 (N393, N317, N349);
xor XOR2_77 (N406, N318, N350);
xor XOR2_78 (N419, N319, N351);
xor XOR2_79 (N432, N320, N352);
xor XOR2_80 (N445, N321, N353);
not NOT1_81 (N554, N354);
not NOT1_82 (N555, N367);
  not NOT1_83 (keyinput_Wire_0[12], N380);
  xor keyGate_0_12(N556, keyinput12, keyinput_Wire_0[12]);
not NOT1_84 (N557, N354);
not NOT1_85 (N558, N367);
not NOT1_86 (N559, N393);
not NOT1_87 (N560, N354);
  not NOT1_88 (keyinput_Wire_0[13], N380);
  xor keyGate_0_13(KeyNOTWire_0[5], keyinput13, keyinput_Wire_0[13]);
  not KeyNOTGate_0_5(N561, KeyNOTWire_0[5]);
not NOT1_89 (N562, N393);
  not NOT1_90 (keyinput_Wire_0[14], N367);
  xnor keyGate_0_14(KeyNOTWire_0[6], keyinput14, keyinput_Wire_0[14]);
  not KeyNOTGate_0_6(N563, KeyNOTWire_0[6]);
not NOT1_91 (N564, N380);
not NOT1_92 (N565, N393);
not NOT1_93 (N566, N419);
  not NOT1_94 (keyinput_Wire_0[15], N445);
  xor keyGate_0_15(N567, keyinput15, keyinput_Wire_0[15]);
not NOT1_95 (N568, N419);
not NOT1_96 (N569, N432);
not NOT1_97 (N570, N406);
not NOT1_98 (N571, N445);
not NOT1_99 (N572, N406);
not NOT1_100 (N573, N432);
not NOT1_101 (N574, N406);
  not NOT1_102 (keyinput_Wire_0[16], N419);
  xor keyGate_0_16(N575, keyinput16, keyinput_Wire_0[16]);
not NOT1_103 (N576, N432);
not NOT1_104 (N577, N406);
not NOT1_105 (N578, N419);
not NOT1_106 (N579, N445);
not NOT1_107 (N580, N406);
not NOT1_108 (N581, N432);
not NOT1_109 (N582, N445);
not NOT1_110 (N583, N419);
not NOT1_111 (N584, N432);
not NOT1_112 (N585, N445);
not NOT1_113 (N586, N367);
not NOT1_114 (N587, N393);
  not NOT1_115 (keyinput_Wire_0[17], N367);
  xor keyGate_0_17(KeyNOTWire_0[7], keyinput17, keyinput_Wire_0[17]);
  not KeyNOTGate_0_7(N588, KeyNOTWire_0[7]);
not NOT1_116 (N589, N380);
  not NOT1_117 (keyinput_Wire_0[18], N354);
  xor keyGate_0_18(N590, keyinput18, keyinput_Wire_0[18]);
  not NOT1_118 (keyinput_Wire_0[19], N393);
  xor keyGate_0_19(KeyNOTWire_0[8], keyinput19, keyinput_Wire_0[19]);
  not KeyNOTGate_0_8(N591, KeyNOTWire_0[8]);
not NOT1_119 (N592, N354);
not NOT1_120 (N593, N380);
and AND4_121 (N594, N554, N555, N556, N393);
and AND4_122 (N595, N557, N558, N380, N559);
and AND4_123 (N596, N560, N367, N561, N562);
and AND4_124 (N597, N354, N563, N564, N565);
  and AND4_125 (keyinput_Wire_0[20], N574, N575, N576, N445);
  xor keyGate_0_20(KeyNOTWire_0[9], keyinput20, keyinput_Wire_0[20]);
  not KeyNOTGate_0_9(N598, KeyNOTWire_0[9]);
and AND4_126 (N599, N577, N578, N432, N579);
and AND4_127 (N600, N580, N419, N581, N582);
and AND4_128 (N601, N406, N583, N584, N585);
or OR4_129 (N602, N594, N595, N596, N597);
or OR4_130 (N607, N598, N599, N600, N601);
and AND5_131 (N620, N406, N566, N432, N567, N602);
and AND5_132 (N625, N406, N568, N569, N445, N602);
and AND5_133 (N630, N570, N419, N432, N571, N602);
and AND5_134 (N635, N572, N419, N573, N445, N602);
and AND5_135 (N640, N354, N586, N380, N587, N607);
and AND5_136 (N645, N354, N588, N589, N393, N607);
and AND5_137 (N650, N590, N367, N380, N591, N607);
and AND5_138 (N655, N592, N367, N593, N393, N607);
  and AND2_139 (keyinput_Wire_0[21], N354, N620);
  xnor keyGate_0_21(KeyNOTWire_0[10], keyinput21, keyinput_Wire_0[21]);
  not KeyNOTGate_0_10(N692, KeyNOTWire_0[10]);
and AND2_140 (N693, N367, N620);
and AND2_141 (N694, N380, N620);
and AND2_142 (N695, N393, N620);
and AND2_143 (N696, N354, N625);
and AND2_144 (N697, N367, N625);
and AND2_145 (N698, N380, N625);
and AND2_146 (N699, N393, N625);
and AND2_147 (N700, N354, N630);
and AND2_148 (N701, N367, N630);
and AND2_149 (N702, N380, N630);
and AND2_150 (N703, N393, N630);
and AND2_151 (N704, N354, N635);
and AND2_152 (N705, N367, N635);
and AND2_153 (N706, N380, N635);
and AND2_154 (N707, N393, N635);
and AND2_155 (N708, N406, N640);
and AND2_156 (N709, N419, N640);
and AND2_157 (N710, N432, N640);
  and AND2_158 (keyinput_Wire_0[22], N445, N640);
  xor keyGate_0_22(KeyNOTWire_0[11], keyinput22, keyinput_Wire_0[22]);
  not KeyNOTGate_0_11(N711, KeyNOTWire_0[11]);
  and AND2_159 (keyinput_Wire_0[23], N406, N645);
  xnor keyGate_0_23(N712, keyinput23, keyinput_Wire_0[23]);
and AND2_160 (N713, N419, N645);
and AND2_161 (N714, N432, N645);
and AND2_162 (N715, N445, N645);
and AND2_163 (N716, N406, N650);
and AND2_164 (N717, N419, N650);
and AND2_165 (N718, N432, N650);
  and AND2_166 (keyinput_Wire_0[24], N445, N650);
  xnor keyGate_0_24(N719, keyinput24, keyinput_Wire_0[24]);
  and AND2_167 (keyinput_Wire_0[25], N406, N655);
  xnor keyGate_0_25(N720, keyinput25, keyinput_Wire_0[25]);
and AND2_168 (N721, N419, N655);
and AND2_169 (N722, N432, N655);
and AND2_170 (N723, N445, N655);
xor XOR2_171 (N724, N1, N692);
xor XOR2_172 (N725, N5, N693);
xor XOR2_173 (N726, N9, N694);
xor XOR2_174 (N727, N13, N695);
xor XOR2_175 (N728, N17, N696);
xor XOR2_176 (N729, N21, N697);
xor XOR2_177 (N730, N25, N698);
  xor XOR2_178 (keyinput_Wire_0[26], N29, N699);
  xor keyGate_0_26(N731, keyinput26, keyinput_Wire_0[26]);
xor XOR2_179 (N732, N33, N700);
xor XOR2_180 (N733, N37, N701);
xor XOR2_181 (N734, N41, N702);
xor XOR2_182 (N735, N45, N703);
xor XOR2_183 (N736, N49, N704);
xor XOR2_184 (N737, N53, N705);
xor XOR2_185 (N738, N57, N706);
xor XOR2_186 (N739, N61, N707);
  xor XOR2_187 (keyinput_Wire_0[27], N65, N708);
  xor keyGate_0_27(KeyNOTWire_0[12], keyinput27, keyinput_Wire_0[27]);
  not KeyNOTGate_0_12(N740, KeyNOTWire_0[12]);
  xor XOR2_188 (keyinput_Wire_0[28], N69, N709);
  xor keyGate_0_28(KeyNOTWire_0[13], keyinput28, keyinput_Wire_0[28]);
  not KeyNOTGate_0_13(N741, KeyNOTWire_0[13]);
xor XOR2_189 (N742, N73, N710);
  xor XOR2_190 (keyinput_Wire_0[29], N77, N711);
  xnor keyGate_0_29(N743, keyinput29, keyinput_Wire_0[29]);
  xor XOR2_191 (keyinput_Wire_0[30], N81, N712);
  xnor keyGate_0_30(KeyNOTWire_0[14], keyinput30, keyinput_Wire_0[30]);
  not KeyNOTGate_0_14(N744, KeyNOTWire_0[14]);
xor XOR2_192 (N745, N85, N713);
  xor XOR2_193 (keyinput_Wire_0[31], N89, N714);
  xor keyGate_0_31(KeyNOTWire_0[15], keyinput31, keyinput_Wire_0[31]);
  not KeyNOTGate_0_15(N746, KeyNOTWire_0[15]);
xor XOR2_194 (N747, N93, N715);
xor XOR2_195 (N748, N97, N716);
xor XOR2_196 (N749, N101, N717);
xor XOR2_197 (N750, N105, N718);
xor XOR2_198 (N751, N109, N719);
xor XOR2_199 (N752, N113, N720);
xor XOR2_200 (KeyWire_0_1, N117, N721);
  xor flip_it (N753, KeyWire_0_1, KeyWire_0_2 );
xor XOR2_201 (N754, N121, N722);
xor XOR2_202 (N755, N125, N723);

AntiSAT some_name( KeyWire_0_2, N57, N130, N135, N132, N41, N136, N17, N49, N137, N13, N125, N85, N77, N29, N81, N61, N89, N21, N133, N9, N53, N121, N113, N109, N73, N65, N129, N131, N69, N5, N45, N33, N101, N37, N25, N93, N117, N1, N134, N97, N105, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
       keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
       keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
       keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
       keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
       keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
       keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
       keyinput144, keyinput145, keyinput146, keyinput147, keyinput148,
       keyinput149, keyinput150, keyinput151, keyinput152, keyinput153,
       keyinput154);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N57, N130, N135, N132, N41, N136, N17, N49, N137, N13, N125, N85, N77, N29, N81, N61, N89, N21, N133, N9, N53, N121, N113, N109, N73, N65, N129, N131, N69, N5, N45, N33, N101, N37, N25, N93, N117, N1, N134, N97, N105, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113 ,
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
        keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
        keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
        keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
        keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
        keyinput144, keyinput145, keyinput146, keyinput147, keyinput148,
        keyinput149, keyinput150, keyinput151, keyinput152, keyinput153,
        keyinput154);

  input keyinput114, keyinput115, keyinput116, keyinput117, keyinput118;
  input keyinput119, keyinput120, keyinput121, keyinput122, keyinput123;
  input keyinput124, keyinput125, keyinput126, keyinput127, keyinput128;
  input keyinput129, keyinput130, keyinput131, keyinput132, keyinput133;
  input keyinput134, keyinput135, keyinput136, keyinput137, keyinput138;
  input keyinput139, keyinput140, keyinput141, keyinput142, keyinput143;
  input keyinput144, keyinput145, keyinput146, keyinput147, keyinput148;
  input keyinput149, keyinput150, keyinput151, keyinput152, keyinput153;
  input keyinput154;

  wire [0:40] keyNTin_Wire_1;
  wire [0:23] KeyNOTWire_1;

  input N57, N130, N135, N132, N41, N136, N17, N49, N137, N13, N125, N85, N77, N29, N81, N61, N89, N21, N133, N9, N53, N121, N113, N109, N73, N65, N129, N131, N69, N5, N45, N33, N101, N37, N25, N93, N117, N1, N134, N97, N105;
  input keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83 ;

  xnor KeyGate0 (keyNTin_Wire_1[0], N57, keyinput32);
  xor keyNTinGate_1_0(newWire_0, keyinput114, keyNTin_Wire_1[0]);
  xor  KeyGate1 (keyNTin_Wire_1[1], N130, keyinput33);
  xor keyNTinGate_1_1(KeyNOTWire_1[0], keyinput115, keyNTin_Wire_1[1]);
  not KeyNOTGate_1_0(newWire_1, KeyNOTWire_1[0]);
  xor  KeyGate2 (keyNTin_Wire_1[2], N135, keyinput34);
  xnor keyNTinGate_1_2(KeyNOTWire_1[1], keyinput116, keyNTin_Wire_1[2]);
  not KeyNOTGate_1_1(newWire_2, KeyNOTWire_1[1]);
  xnor KeyGate3 (keyNTin_Wire_1[3], N132, keyinput35);
  xnor keyNTinGate_1_3(KeyNOTWire_1[2], keyinput117, keyNTin_Wire_1[3]);
  not KeyNOTGate_1_2(newWire_3, KeyNOTWire_1[2]);
  xor  KeyGate4 (keyNTin_Wire_1[4], N41, keyinput36);
  xor keyNTinGate_1_4(newWire_4, keyinput118, keyNTin_Wire_1[4]);
  xnor KeyGate5 (keyNTin_Wire_1[5], N136, keyinput37);
  xnor keyNTinGate_1_5(newWire_5, keyinput119, keyNTin_Wire_1[5]);
  xnor KeyGate6 (keyNTin_Wire_1[6], N17, keyinput38);
  xor keyNTinGate_1_6(KeyNOTWire_1[3], keyinput120, keyNTin_Wire_1[6]);
  not KeyNOTGate_1_3(newWire_6, KeyNOTWire_1[3]);
  xnor KeyGate7 (keyNTin_Wire_1[7], N49, keyinput39);
  xnor keyNTinGate_1_7(KeyNOTWire_1[4], keyinput121, keyNTin_Wire_1[7]);
  not KeyNOTGate_1_4(newWire_7, KeyNOTWire_1[4]);
  xor  KeyGate8 (keyNTin_Wire_1[8], N137, keyinput40);
  xor keyNTinGate_1_8(newWire_8, keyinput122, keyNTin_Wire_1[8]);
  xnor KeyGate9 (newWire_9, N13, keyinput41);
  xnor KeyGate10 (newWire_10, N125, keyinput42);
  xnor KeyGate11 (keyNTin_Wire_1[9], N85, keyinput43);
  xnor keyNTinGate_1_9(KeyNOTWire_1[5], keyinput123, keyNTin_Wire_1[9]);
  not KeyNOTGate_1_5(newWire_11, KeyNOTWire_1[5]);
  xnor KeyGate12 (keyNTin_Wire_1[10], N77, keyinput44);
  xnor keyNTinGate_1_10(KeyNOTWire_1[6], keyinput124, keyNTin_Wire_1[10]);
  not KeyNOTGate_1_6(newWire_12, KeyNOTWire_1[6]);
  xnor KeyGate13 (newWire_13, N29, keyinput45);
  xor  KeyGate14 (keyNTin_Wire_1[11], N81, keyinput46);
  xnor keyNTinGate_1_11(KeyNOTWire_1[7], keyinput125, keyNTin_Wire_1[11]);
  not KeyNOTGate_1_7(newWire_14, KeyNOTWire_1[7]);
  xnor KeyGate15 (keyNTin_Wire_1[12], N61, keyinput47);
  xor keyNTinGate_1_12(KeyNOTWire_1[8], keyinput126, keyNTin_Wire_1[12]);
  not KeyNOTGate_1_8(newWire_15, KeyNOTWire_1[8]);
  xnor KeyGate16 (keyNTin_Wire_1[13], N89, keyinput48);
  xnor keyNTinGate_1_13(newWire_16, keyinput127, keyNTin_Wire_1[13]);
  xnor KeyGate17 (newWire_17, N21, keyinput49);
  xnor KeyGate18 (newWire_18, N133, keyinput50);
  xnor KeyGate19 (newWire_19, N9, keyinput51);
  xnor KeyGate20 (newWire_20, N53, keyinput52);
  xor  KeyGate21 (keyNTin_Wire_1[14], N121, keyinput53);
  xor keyNTinGate_1_14(KeyNOTWire_1[9], keyinput128, keyNTin_Wire_1[14]);
  not KeyNOTGate_1_9(newWire_21, KeyNOTWire_1[9]);
  xor  KeyGate22 (newWire_22, N113, keyinput54);
  xor  KeyGate23 (newWire_23, N109, keyinput55);
  xnor KeyGate24 (newWire_24, N73, keyinput56);
  xor  KeyGate25 (newWire_25, N65, keyinput57);
  xnor KeyGate26 (newWire_26, N129, keyinput58);
  xor  KeyGate27 (keyNTin_Wire_1[15], N131, keyinput59);
  xor keyNTinGate_1_15(newWire_27, keyinput129, keyNTin_Wire_1[15]);
  xor  KeyGate28 (keyNTin_Wire_1[16], N69, keyinput60);
  xnor keyNTinGate_1_16(newWire_28, keyinput130, keyNTin_Wire_1[16]);
  xor  KeyGate29 (keyNTin_Wire_1[17], N5, keyinput61);
  xnor keyNTinGate_1_17(KeyNOTWire_1[10], keyinput131, keyNTin_Wire_1[17]);
  not KeyNOTGate_1_10(newWire_29, KeyNOTWire_1[10]);
  xnor KeyGate30 (keyNTin_Wire_1[18], N45, keyinput62);
  xor keyNTinGate_1_18(KeyNOTWire_1[11], keyinput132, keyNTin_Wire_1[18]);
  not KeyNOTGate_1_11(newWire_30, KeyNOTWire_1[11]);
  xor  KeyGate31 (newWire_31, N33, keyinput63);
  xnor KeyGate32 (keyNTin_Wire_1[19], N101, keyinput64);
  xnor keyNTinGate_1_19(KeyNOTWire_1[12], keyinput133, keyNTin_Wire_1[19]);
  not KeyNOTGate_1_12(newWire_32, KeyNOTWire_1[12]);
  xor  KeyGate33 (newWire_33, N37, keyinput65);
  xor  KeyGate34 (keyNTin_Wire_1[20], N25, keyinput66);
  xor keyNTinGate_1_20(KeyNOTWire_1[13], keyinput134, keyNTin_Wire_1[20]);
  not KeyNOTGate_1_13(newWire_34, KeyNOTWire_1[13]);
  xor  KeyGate35 (keyNTin_Wire_1[21], N93, keyinput67);
  xnor keyNTinGate_1_21(newWire_35, keyinput135, keyNTin_Wire_1[21]);
  xor  KeyGate36 (newWire_36, N117, keyinput68);
  xnor KeyGate37 (newWire_37, N1, keyinput69);
  xor  KeyGate38 (newWire_38, N134, keyinput70);
  xor  KeyGate39 (keyNTin_Wire_1[22], N97, keyinput71);
  xor keyNTinGate_1_22(newWire_39, keyinput136, keyNTin_Wire_1[22]);
  xor  KeyGate40 (keyNTin_Wire_1[23], N105, keyinput72);
  xnor keyNTinGate_1_23(newWire_40, keyinput137, keyNTin_Wire_1[23]);
  xor  KeyGate41 (newWire_41, N57, keyinput73);
  xor  KeyGate42 (keyNTin_Wire_1[24], N130, keyinput74);
  xnor keyNTinGate_1_24(newWire_42, keyinput138, keyNTin_Wire_1[24]);
  xor  KeyGate43 (newWire_43, N135, keyinput75);
  xor  KeyGate44 (keyNTin_Wire_1[25], N132, keyinput76);
  xor keyNTinGate_1_25(newWire_44, keyinput139, keyNTin_Wire_1[25]);
  xor  KeyGate45 (newWire_45, N41, keyinput77);
  xor  KeyGate46 (newWire_46, N136, keyinput78);
  xor  KeyGate47 (newWire_47, N17, keyinput79);
  xnor KeyGate48 (keyNTin_Wire_1[26], N49, keyinput80);
  xor keyNTinGate_1_26(KeyNOTWire_1[14], keyinput140, keyNTin_Wire_1[26]);
  not KeyNOTGate_1_14(newWire_48, KeyNOTWire_1[14]);
  xor  KeyGate49 (keyNTin_Wire_1[27], N137, keyinput81);
  xor keyNTinGate_1_27(newWire_49, keyinput141, keyNTin_Wire_1[27]);
  xor  KeyGate50 (keyNTin_Wire_1[28], N13, keyinput82);
  xnor keyNTinGate_1_28(KeyNOTWire_1[15], keyinput142, keyNTin_Wire_1[28]);
  not KeyNOTGate_1_15(newWire_50, KeyNOTWire_1[15]);
  xnor KeyGate51 (keyNTin_Wire_1[29], N125, keyinput83);
  xnor keyNTinGate_1_29(KeyNOTWire_1[16], keyinput143, keyNTin_Wire_1[29]);
  not KeyNOTGate_1_16(newWire_51, KeyNOTWire_1[16]);
  xor  KeyGate52 (keyNTin_Wire_1[30], N85, keyinput84);
  xor keyNTinGate_1_30(KeyNOTWire_1[17], keyinput144, keyNTin_Wire_1[30]);
  not KeyNOTGate_1_17(newWire_52, KeyNOTWire_1[17]);
  xnor KeyGate53 (newWire_53, N77, keyinput85);
  xnor KeyGate54 (newWire_54, N29, keyinput86);
  xnor KeyGate55 (newWire_55, N81, keyinput87);
  xor  KeyGate56 (keyNTin_Wire_1[31], N61, keyinput88);
  xor keyNTinGate_1_31(KeyNOTWire_1[18], keyinput145, keyNTin_Wire_1[31]);
  not KeyNOTGate_1_18(newWire_56, KeyNOTWire_1[18]);
  xnor KeyGate57 (keyNTin_Wire_1[32], N89, keyinput89);
  xnor keyNTinGate_1_32(newWire_57, keyinput146, keyNTin_Wire_1[32]);
  xor  KeyGate58 (newWire_58, N21, keyinput90);
  xor  KeyGate59 (newWire_59, N133, keyinput91);
  xor  KeyGate60 (newWire_60, N9, keyinput92);
  xor  KeyGate61 (newWire_61, N53, keyinput93);
  xnor KeyGate62 (newWire_62, N121, keyinput94);
  xnor KeyGate63 (newWire_63, N113, keyinput95);
  xnor KeyGate64 (keyNTin_Wire_1[33], N109, keyinput96);
  xor keyNTinGate_1_33(newWire_64, keyinput147, keyNTin_Wire_1[33]);
  xnor KeyGate65 (keyNTin_Wire_1[34], N73, keyinput97);
  xnor keyNTinGate_1_34(KeyNOTWire_1[19], keyinput148, keyNTin_Wire_1[34]);
  not KeyNOTGate_1_19(newWire_65, KeyNOTWire_1[19]);
  xnor KeyGate66 (newWire_66, N65, keyinput98);
  xor  KeyGate67 (newWire_67, N129, keyinput99);
  xnor KeyGate68 (newWire_68, N131, keyinput100);
  xor  KeyGate69 (keyNTin_Wire_1[35], N69, keyinput101);
  xor keyNTinGate_1_35(KeyNOTWire_1[20], keyinput149, keyNTin_Wire_1[35]);
  not KeyNOTGate_1_20(newWire_69, KeyNOTWire_1[20]);
  xnor KeyGate70 (newWire_70, N5, keyinput102);
  xor  KeyGate71 (keyNTin_Wire_1[36], N45, keyinput103);
  xnor keyNTinGate_1_36(newWire_71, keyinput150, keyNTin_Wire_1[36]);
  xnor KeyGate72 (newWire_72, N33, keyinput104);
  xnor KeyGate73 (keyNTin_Wire_1[37], N101, keyinput105);
  xnor keyNTinGate_1_37(KeyNOTWire_1[21], keyinput151, keyNTin_Wire_1[37]);
  not KeyNOTGate_1_21(newWire_73, KeyNOTWire_1[21]);
  xor  KeyGate74 (newWire_74, N37, keyinput106);
  xor  KeyGate75 (newWire_75, N25, keyinput107);
  xnor KeyGate76 (newWire_76, N93, keyinput108);
  xor  KeyGate77 (newWire_77, N117, keyinput109);
  xor  KeyGate78 (keyNTin_Wire_1[38], N1, keyinput110);
  xor keyNTinGate_1_38(KeyNOTWire_1[22], keyinput152, keyNTin_Wire_1[38]);
  not KeyNOTGate_1_22(newWire_78, KeyNOTWire_1[22]);
  xnor KeyGate79 (keyNTin_Wire_1[39], N134, keyinput111);
  xnor keyNTinGate_1_39(newWire_79, keyinput153, keyNTin_Wire_1[39]);
  xnor KeyGate80 (newWire_80, N97, keyinput112);
  xnor KeyGate81 (keyNTin_Wire_1[40], N105, keyinput113);
  xor keyNTinGate_1_40(KeyNOTWire_1[23], keyinput154, keyNTin_Wire_1[40]);
  not KeyNOTGate_1_23(newWire_81, KeyNOTWire_1[23]);
  and some_function (newWire_82, newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40 );
  nand compl_function (newWire_83, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81);
  and finalAND (KeyWire_0_2, newWire_82, newWire_83);

endmodule /* AntiSAT */
