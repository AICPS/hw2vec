`timescale 1ns / 1ps
// Verilog
// c432
// Ninputs 36
// Noutputs 7
// NtotalGates 160
// NOT1 40
// NAND2 64
// NOR2 19
// AND9 3
// XOR2 18
// NAND4 14
// AND8 1
// NAND3 1

module top (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
                  N430,N431,N432,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
                  keyinput30, keyinput31,
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36,
        keyinput37, keyinput38, keyinput39, keyinput40, keyinput41,
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46,
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51,
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56,
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61,
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66,
        keyinput67, keyinput68, keyinput69, keyinput70, keyinput71,
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76,
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81,
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86,
        keyinput87, keyinput88, keyinput89, keyinput90, keyinput91,
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96,
        keyinput97, keyinput98, keyinput99, keyinput100, keyinput101,
                  keyinput102, keyinput103,
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
        keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
        keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
        keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
        keyinput139);

  input keyinput104, keyinput105, keyinput106, keyinput107, keyinput108;
  input keyinput109, keyinput110, keyinput111, keyinput112, keyinput113;
  input keyinput114, keyinput115, keyinput116, keyinput117, keyinput118;
  input keyinput119, keyinput120, keyinput121, keyinput122, keyinput123;
  input keyinput124, keyinput125, keyinput126, keyinput127, keyinput128;
  input keyinput129, keyinput130, keyinput131, keyinput132, keyinput133;
  input keyinput134, keyinput135, keyinput136, keyinput137, keyinput138;
  input keyinput139;


  input keyinput32, keyinput33, keyinput34, keyinput35, keyinput36;
  input keyinput37, keyinput38, keyinput39, keyinput40, keyinput41;
  input keyinput42, keyinput43, keyinput44, keyinput45, keyinput46;
  input keyinput47, keyinput48, keyinput49, keyinput50, keyinput51;
  input keyinput52, keyinput53, keyinput54, keyinput55, keyinput56;
  input keyinput57, keyinput58, keyinput59, keyinput60, keyinput61;
  input keyinput62, keyinput63, keyinput64, keyinput65, keyinput66;
  input keyinput67, keyinput68, keyinput69, keyinput70, keyinput71;
  input keyinput72, keyinput73, keyinput74, keyinput75, keyinput76;
  input keyinput77, keyinput78, keyinput79, keyinput80, keyinput81;
  input keyinput82, keyinput83, keyinput84, keyinput85, keyinput86;
  input keyinput87, keyinput88, keyinput89, keyinput90, keyinput91;
  input keyinput92, keyinput93, keyinput94, keyinput95, keyinput96;
  input keyinput97, keyinput98, keyinput99, keyinput100, keyinput101;
  input keyinput102, keyinput103;

  wire KeyWire_0_1 , KeyWire_0_2;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31;

  wire [0:31] keyinput_Wire_0;
  wire [0:17] KeyNOTWire_0;

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;

output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429;

  not NOT1_1 (keyinput_Wire_0[0], N1);
  xnor keyGate_0_0(N118, keyinput0, keyinput_Wire_0[0]);
not NOT1_2 (N119, N4);
  not NOT1_3 (keyinput_Wire_0[1], N11);
  xor keyGate_0_1(N122, keyinput1, keyinput_Wire_0[1]);
not NOT1_4 (N123, N17);
  not NOT1_5 (keyinput_Wire_0[2], N24);
  xnor keyGate_0_2(N126, keyinput2, keyinput_Wire_0[2]);
  not NOT1_6 (keyinput_Wire_0[3], N30);
  xnor keyGate_0_3(N127, keyinput3, keyinput_Wire_0[3]);
  not NOT1_7 (keyinput_Wire_0[4], N37);
  xor keyGate_0_4(KeyNOTWire_0[0], keyinput4, keyinput_Wire_0[4]);
  not KeyNOTGate_0_0(N130, KeyNOTWire_0[0]);
not NOT1_8 (N131, N43);
  not NOT1_9 (keyinput_Wire_0[5], N50);
  xnor keyGate_0_5(KeyNOTWire_0[1], keyinput5, keyinput_Wire_0[5]);
  not KeyNOTGate_0_1(N134, KeyNOTWire_0[1]);
not NOT1_10 (N135, N56);
  not NOT1_11 (keyinput_Wire_0[6], N63);
  xor keyGate_0_6(KeyNOTWire_0[2], keyinput6, keyinput_Wire_0[6]);
  not KeyNOTGate_0_2(N138, KeyNOTWire_0[2]);
not NOT1_12 (N139, N69);
  not NOT1_13 (keyinput_Wire_0[7], N76);
  xnor keyGate_0_7(KeyNOTWire_0[3], keyinput7, keyinput_Wire_0[7]);
  not KeyNOTGate_0_3(N142, KeyNOTWire_0[3]);
not NOT1_14 (N143, N82);
  not NOT1_15 (keyinput_Wire_0[8], N89);
  xnor keyGate_0_8(KeyNOTWire_0[4], keyinput8, keyinput_Wire_0[8]);
  not KeyNOTGate_0_4(N146, KeyNOTWire_0[4]);
  not NOT1_16 (keyinput_Wire_0[9], N95);
  xnor keyGate_0_9(KeyNOTWire_0[5], keyinput9, keyinput_Wire_0[9]);
  not KeyNOTGate_0_5(N147, KeyNOTWire_0[5]);
  not NOT1_17 (keyinput_Wire_0[10], N102);
  xnor keyGate_0_10(KeyNOTWire_0[6], keyinput10, keyinput_Wire_0[10]);
  not KeyNOTGate_0_6(N150, KeyNOTWire_0[6]);
not NOT1_18 (N151, N108);
  nand NAND2_19 (keyinput_Wire_0[11], N118, N4);
  xnor keyGate_0_11(N154, keyinput11, keyinput_Wire_0[11]);
nor NOR2_20 (N157, N8, N119);
nor NOR2_21 (N158, N14, N119);
  nand NAND2_22 (keyinput_Wire_0[12], N122, N17);
  xor keyGate_0_12(KeyNOTWire_0[7], keyinput12, keyinput_Wire_0[12]);
  not KeyNOTGate_0_7(N159, KeyNOTWire_0[7]);
  nand NAND2_23 (keyinput_Wire_0[13], N126, N30);
  xnor keyGate_0_13(KeyNOTWire_0[8], keyinput13, keyinput_Wire_0[13]);
  not KeyNOTGate_0_8(N162, KeyNOTWire_0[8]);
  nand NAND2_24 (keyinput_Wire_0[14], N130, N43);
  xor keyGate_0_14(KeyNOTWire_0[9], keyinput14, keyinput_Wire_0[14]);
  not KeyNOTGate_0_9(N165, KeyNOTWire_0[9]);
  nand NAND2_25 (keyinput_Wire_0[15], N134, N56);
  xor keyGate_0_15(KeyNOTWire_0[10], keyinput15, keyinput_Wire_0[15]);
  not KeyNOTGate_0_10(N168, KeyNOTWire_0[10]);
  nand NAND2_26 (keyinput_Wire_0[16], N138, N69);
  xnor keyGate_0_16(N171, keyinput16, keyinput_Wire_0[16]);
  nand NAND2_27 (keyinput_Wire_0[17], N142, N82);
  xor keyGate_0_17(N174, keyinput17, keyinput_Wire_0[17]);
  nand NAND2_28 (keyinput_Wire_0[18], N146, N95);
  xor keyGate_0_18(KeyNOTWire_0[11], keyinput18, keyinput_Wire_0[18]);
  not KeyNOTGate_0_11(N177, KeyNOTWire_0[11]);
  nand NAND2_29 (keyinput_Wire_0[19], N150, N108);
  xor keyGate_0_19(N180, keyinput19, keyinput_Wire_0[19]);
nor NOR2_30 (N183, N21, N123);
nor NOR2_31 (N184, N27, N123);
nor NOR2_32 (N185, N34, N127);
  nor NOR2_33 (keyinput_Wire_0[20], N40, N127);
  xnor keyGate_0_20(KeyNOTWire_0[12], keyinput20, keyinput_Wire_0[20]);
  not KeyNOTGate_0_12(N186, KeyNOTWire_0[12]);
nor NOR2_34 (N187, N47, N131);
nor NOR2_35 (N188, N53, N131);
nor NOR2_36 (N189, N60, N135);
nor NOR2_37 (N190, N66, N135);
nor NOR2_38 (N191, N73, N139);
nor NOR2_39 (N192, N79, N139);
nor NOR2_40 (N193, N86, N143);
nor NOR2_41 (N194, N92, N143);
nor NOR2_42 (N195, N99, N147);
  nor NOR2_43 (keyinput_Wire_0[21], N105, N147);
  xor keyGate_0_21(N196, keyinput21, keyinput_Wire_0[21]);
nor NOR2_44 (N197, N112, N151);
nor NOR2_45 (N198, N115, N151);
  and AND9_46 (keyinput_Wire_0[22], N154, N159, N162, N165, N168, N171, N174, N177, N180);
  xnor keyGate_0_22(N199, keyinput22, keyinput_Wire_0[22]);
  not NOT1_47 (keyinput_Wire_0[23], N199);
  xnor keyGate_0_23(KeyNOTWire_0[13], keyinput23, keyinput_Wire_0[23]);
  not KeyNOTGate_0_13(N203, KeyNOTWire_0[13]);
not NOT1_48 (N213, N199);
not NOT1_49 (N223, N199);
xor XOR2_50 (N224, N203, N154);
xor XOR2_51 (N227, N203, N159);
  xor XOR2_52 (keyinput_Wire_0[24], N203, N162);
  xor keyGate_0_24(KeyNOTWire_0[14], keyinput24, keyinput_Wire_0[24]);
  not KeyNOTGate_0_14(N230, KeyNOTWire_0[14]);
  xor XOR2_53 (keyinput_Wire_0[25], N203, N165);
  xnor keyGate_0_25(N233, keyinput25, keyinput_Wire_0[25]);
xor XOR2_54 (N236, N203, N168);
xor XOR2_55 (N239, N203, N171);
nand NAND2_56 (N242, N1, N213);
xor XOR2_57 (N243, N203, N174);
nand NAND2_58 (N246, N213, N11);
xor XOR2_59 (N247, N203, N177);
nand NAND2_60 (N250, N213, N24);
xor XOR2_61 (N251, N203, N180);
nand NAND2_62 (N254, N213, N37);
nand NAND2_63 (N255, N213, N50);
nand NAND2_64 (N256, N213, N63);
nand NAND2_65 (N257, N213, N76);
nand NAND2_66 (N258, N213, N89);
nand NAND2_67 (N259, N213, N102);
nand NAND2_68 (N260, N224, N157);
nand NAND2_69 (N263, N224, N158);
nand NAND2_70 (N264, N227, N183);
nand NAND2_71 (N267, N230, N185);
nand NAND2_72 (N270, N233, N187);
nand NAND2_73 (N273, N236, N189);
nand NAND2_74 (N276, N239, N191);
nand NAND2_75 (N279, N243, N193);
nand NAND2_76 (N282, N247, N195);
nand NAND2_77 (N285, N251, N197);
nand NAND2_78 (N288, N227, N184);
  nand NAND2_79 (keyinput_Wire_0[26], N230, N186);
  xnor keyGate_0_26(N289, keyinput26, keyinput_Wire_0[26]);
nand NAND2_80 (N290, N233, N188);
nand NAND2_81 (N291, N236, N190);
nand NAND2_82 (N292, N239, N192);
nand NAND2_83 (N293, N243, N194);
nand NAND2_84 (N294, N247, N196);
nand NAND2_85 (N295, N251, N198);
and AND9_86 (N296, N260, N264, N267, N270, N273, N276, N279, N282, N285);
not NOT1_87 (N300, N263);
not NOT1_88 (N301, N288);
  not NOT1_89 (keyinput_Wire_0[27], N289);
  xnor keyGate_0_27(N302, keyinput27, keyinput_Wire_0[27]);
  not NOT1_90 (keyinput_Wire_0[28], N290);
  xnor keyGate_0_28(KeyNOTWire_0[15], keyinput28, keyinput_Wire_0[28]);
  not KeyNOTGate_0_15(N303, KeyNOTWire_0[15]);
not NOT1_91 (N304, N291);
not NOT1_92 (N305, N292);
not NOT1_93 (N306, N293);
not NOT1_94 (N307, N294);
not NOT1_95 (N308, N295);
not NOT1_96 (N309, N296);
not NOT1_97 (N319, N296);
not NOT1_98 (N329, N296);
xor XOR2_99 (N330, N309, N260);
xor XOR2_100 (N331, N309, N264);
xor XOR2_101 (N332, N309, N267);
xor XOR2_102 (N333, N309, N270);
nand NAND2_103 (N334, N8, N319);
xor XOR2_104 (N335, N309, N273);
nand NAND2_105 (N336, N319, N21);
xor XOR2_106 (N337, N309, N276);
nand NAND2_107 (N338, N319, N34);
  xor XOR2_108 (keyinput_Wire_0[29], N309, N279);
  xnor keyGate_0_29(KeyNOTWire_0[16], keyinput29, keyinput_Wire_0[29]);
  not KeyNOTGate_0_16(N339, KeyNOTWire_0[16]);
nand NAND2_109 (N340, N319, N47);
xor XOR2_110 (N341, N309, N282);
nand NAND2_111 (N342, N319, N60);
xor XOR2_112 (N343, N309, N285);
nand NAND2_113 (N344, N319, N73);
nand NAND2_114 (N345, N319, N86);
nand NAND2_115 (N346, N319, N99);
nand NAND2_116 (N347, N319, N112);
nand NAND2_117 (N348, N330, N300);
nand NAND2_118 (N349, N331, N301);
nand NAND2_119 (N350, N332, N302);
nand NAND2_120 (N351, N333, N303);
nand NAND2_121 (N352, N335, N304);
nand NAND2_122 (N353, N337, N305);
nand NAND2_123 (N354, N339, N306);
nand NAND2_124 (N355, N341, N307);
nand NAND2_125 (N356, N343, N308);
and AND9_126 (N357, N348, N349, N350, N351, N352, N353, N354, N355, N356);
  not NOT1_127 (keyinput_Wire_0[30], N357);
  xor keyGate_0_30(KeyNOTWire_0[17], keyinput30, keyinput_Wire_0[30]);
  not KeyNOTGate_0_17(N360, KeyNOTWire_0[17]);
not NOT1_128 (N370, N357);
nand NAND2_129 (N371, N14, N360);
nand NAND2_130 (N372, N360, N27);
nand NAND2_131 (N373, N360, N40);
nand NAND2_132 (N374, N360, N53);
nand NAND2_133 (N375, N360, N66);
nand NAND2_134 (N376, N360, N79);
nand NAND2_135 (N377, N360, N92);
  nand NAND2_136 (keyinput_Wire_0[31], N360, N105);
  xor keyGate_0_31(N378, keyinput31, keyinput_Wire_0[31]);
nand NAND2_137 (N379, N360, N115);
nand NAND4_138 (N380, N4, N242, N334, N371);
nand NAND4_139 (N381, N246, N336, N372, N17);
nand NAND4_140 (N386, N250, N338, N373, N30);
nand NAND4_141 (N393, N254, N340, N374, N43);
nand NAND4_142 (N399, N255, N342, N375, N56);
nand NAND4_143 (N404, N256, N344, N376, N69);
nand NAND4_144 (N407, N257, N345, N377, N82);
nand NAND4_145 (N411, N258, N346, N378, N95);
nand NAND4_146 (N414, N259, N347, N379, N108);
not NOT1_147 (N415, N380);
and AND8_148 (N416, N381, N386, N393, N399, N404, N407, N411, N414);
not NOT1_149 (N417, N393);
not NOT1_150 (N418, N404);
not NOT1_151 (N419, N407);
not NOT1_152 (N420, N411);
nor NOR2_153 (N421, N415, N416);
nand NAND2_154 (N422, N386, N417);
nand NAND4_155 (N425, N386, N393, N418, N399);
nand NAND3_156 (N428, N399, N393, N419);
nand NAND4_157 (N429, N386, N393, N407, N420);
nand NAND4_158 (N430, N381, N386, N422, N399);
nand NAND4_159 (KeyWire_0_1, N381, N386, N425, N428);
  xor flip_it (N431, KeyWire_0_1, KeyWire_0_2 );
nand NAND4_160 (N432, N381, N422, N425, N429);

AntiSAT some_name( KeyWire_0_2, N60, N37, N53, N4, N69, N1, N43, N99, N34, N112, N30, N21, N8, N24, N17, N102, N47, N56, N79, N40, N73, N89, N95, N11, N27, N115, N66, N50, N92, N86, N63, N82, N105, N76, N108, N14, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
       keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
       keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
       keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
       keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
       keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
       keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
       keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
       keyinput139);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N60, N37, N53, N4, N69, N1, N43, N99, N34, N112, N30, N21, N8, N24, N17, N102, N47, N56, N79, N40, N73, N89, N95, N11, N27, N115, N66, N50, N92, N86, N63, N82, N105, N76, N108, N14, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103 ,
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
        keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
        keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
        keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
        keyinput139);

  input keyinput104, keyinput105, keyinput106, keyinput107, keyinput108;
  input keyinput109, keyinput110, keyinput111, keyinput112, keyinput113;
  input keyinput114, keyinput115, keyinput116, keyinput117, keyinput118;
  input keyinput119, keyinput120, keyinput121, keyinput122, keyinput123;
  input keyinput124, keyinput125, keyinput126, keyinput127, keyinput128;
  input keyinput129, keyinput130, keyinput131, keyinput132, keyinput133;
  input keyinput134, keyinput135, keyinput136, keyinput137, keyinput138;
  input keyinput139;

  wire [0:35] keyNTin_Wire_1;
  wire [0:19] KeyNOTWire_1;

  input N60, N37, N53, N4, N69, N1, N43, N99, N34, N112, N30, N21, N8, N24, N17, N102, N47, N56, N79, N40, N73, N89, N95, N11, N27, N115, N66, N50, N92, N86, N63, N82, N105, N76, N108, N14;
  input keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73 ;

  xor  KeyGate0 (newWire_0, N60, keyinput32);
  xor  KeyGate1 (newWire_1, N37, keyinput33);
  xnor KeyGate2 (newWire_2, N53, keyinput34);
  xor  KeyGate3 (keyNTin_Wire_1[0], N4, keyinput35);
  xnor keyNTinGate_1_0(KeyNOTWire_1[0], keyinput104, keyNTin_Wire_1[0]);
  not KeyNOTGate_1_0(newWire_3, KeyNOTWire_1[0]);
  xor  KeyGate4 (newWire_4, N69, keyinput36);
  xnor KeyGate5 (newWire_5, N1, keyinput37);
  xor  KeyGate6 (keyNTin_Wire_1[1], N43, keyinput38);
  xor keyNTinGate_1_1(newWire_6, keyinput105, keyNTin_Wire_1[1]);
  xnor KeyGate7 (keyNTin_Wire_1[2], N99, keyinput39);
  xor keyNTinGate_1_2(newWire_7, keyinput106, keyNTin_Wire_1[2]);
  xnor KeyGate8 (keyNTin_Wire_1[3], N34, keyinput40);
  xor keyNTinGate_1_3(KeyNOTWire_1[1], keyinput107, keyNTin_Wire_1[3]);
  not KeyNOTGate_1_1(newWire_8, KeyNOTWire_1[1]);
  xnor KeyGate9 (keyNTin_Wire_1[4], N112, keyinput41);
  xnor keyNTinGate_1_4(KeyNOTWire_1[2], keyinput108, keyNTin_Wire_1[4]);
  not KeyNOTGate_1_2(newWire_9, KeyNOTWire_1[2]);
  xnor KeyGate10 (keyNTin_Wire_1[5], N30, keyinput42);
  xnor keyNTinGate_1_5(newWire_10, keyinput109, keyNTin_Wire_1[5]);
  xor  KeyGate11 (newWire_11, N21, keyinput43);
  xnor KeyGate12 (newWire_12, N8, keyinput44);
  xor  KeyGate13 (keyNTin_Wire_1[6], N24, keyinput45);
  xnor keyNTinGate_1_6(newWire_13, keyinput110, keyNTin_Wire_1[6]);
  xnor KeyGate14 (newWire_14, N17, keyinput46);
  xnor KeyGate15 (newWire_15, N102, keyinput47);
  xnor KeyGate16 (keyNTin_Wire_1[7], N47, keyinput48);
  xnor keyNTinGate_1_7(KeyNOTWire_1[3], keyinput111, keyNTin_Wire_1[7]);
  not KeyNOTGate_1_3(newWire_16, KeyNOTWire_1[3]);
  xor  KeyGate17 (keyNTin_Wire_1[8], N56, keyinput49);
  xnor keyNTinGate_1_8(KeyNOTWire_1[4], keyinput112, keyNTin_Wire_1[8]);
  not KeyNOTGate_1_4(newWire_17, KeyNOTWire_1[4]);
  xnor KeyGate18 (keyNTin_Wire_1[9], N79, keyinput50);
  xnor keyNTinGate_1_9(newWire_18, keyinput113, keyNTin_Wire_1[9]);
  xnor KeyGate19 (keyNTin_Wire_1[10], N40, keyinput51);
  xor keyNTinGate_1_10(newWire_19, keyinput114, keyNTin_Wire_1[10]);
  xor  KeyGate20 (newWire_20, N73, keyinput52);
  xor  KeyGate21 (keyNTin_Wire_1[11], N89, keyinput53);
  xnor keyNTinGate_1_11(newWire_21, keyinput115, keyNTin_Wire_1[11]);
  xor  KeyGate22 (newWire_22, N95, keyinput54);
  xor  KeyGate23 (keyNTin_Wire_1[12], N11, keyinput55);
  xnor keyNTinGate_1_12(KeyNOTWire_1[5], keyinput116, keyNTin_Wire_1[12]);
  not KeyNOTGate_1_5(newWire_23, KeyNOTWire_1[5]);
  xor  KeyGate24 (keyNTin_Wire_1[13], N27, keyinput56);
  xor keyNTinGate_1_13(KeyNOTWire_1[6], keyinput117, keyNTin_Wire_1[13]);
  not KeyNOTGate_1_6(newWire_24, KeyNOTWire_1[6]);
  xor  KeyGate25 (keyNTin_Wire_1[14], N115, keyinput57);
  xor keyNTinGate_1_14(newWire_25, keyinput118, keyNTin_Wire_1[14]);
  xor  KeyGate26 (keyNTin_Wire_1[15], N66, keyinput58);
  xnor keyNTinGate_1_15(newWire_26, keyinput119, keyNTin_Wire_1[15]);
  xnor KeyGate27 (keyNTin_Wire_1[16], N50, keyinput59);
  xnor keyNTinGate_1_16(KeyNOTWire_1[7], keyinput120, keyNTin_Wire_1[16]);
  not KeyNOTGate_1_7(newWire_27, KeyNOTWire_1[7]);
  xnor KeyGate28 (keyNTin_Wire_1[17], N92, keyinput60);
  xor keyNTinGate_1_17(KeyNOTWire_1[8], keyinput121, keyNTin_Wire_1[17]);
  not KeyNOTGate_1_8(newWire_28, KeyNOTWire_1[8]);
  xnor KeyGate29 (keyNTin_Wire_1[18], N86, keyinput61);
  xor keyNTinGate_1_18(KeyNOTWire_1[9], keyinput122, keyNTin_Wire_1[18]);
  not KeyNOTGate_1_9(newWire_29, KeyNOTWire_1[9]);
  xor  KeyGate30 (newWire_30, N63, keyinput62);
  xor  KeyGate31 (keyNTin_Wire_1[19], N82, keyinput63);
  xor keyNTinGate_1_19(KeyNOTWire_1[10], keyinput123, keyNTin_Wire_1[19]);
  not KeyNOTGate_1_10(newWire_31, KeyNOTWire_1[10]);
  xnor KeyGate32 (keyNTin_Wire_1[20], N105, keyinput64);
  xor keyNTinGate_1_20(KeyNOTWire_1[11], keyinput124, keyNTin_Wire_1[20]);
  not KeyNOTGate_1_11(newWire_32, KeyNOTWire_1[11]);
  xor  KeyGate33 (keyNTin_Wire_1[21], N76, keyinput65);
  xor keyNTinGate_1_21(newWire_33, keyinput125, keyNTin_Wire_1[21]);
  xnor KeyGate34 (newWire_34, N108, keyinput66);
  xor  KeyGate35 (newWire_35, N14, keyinput67);
  xor  KeyGate36 (newWire_36, N60, keyinput68);
  xnor KeyGate37 (keyNTin_Wire_1[22], N37, keyinput69);
  xor keyNTinGate_1_22(newWire_37, keyinput126, keyNTin_Wire_1[22]);
  xnor KeyGate38 (newWire_38, N53, keyinput70);
  xor  KeyGate39 (newWire_39, N4, keyinput71);
  xor  KeyGate40 (keyNTin_Wire_1[23], N69, keyinput72);
  xor keyNTinGate_1_23(newWire_40, keyinput127, keyNTin_Wire_1[23]);
  xnor KeyGate41 (newWire_41, N1, keyinput73);
  xor  KeyGate42 (newWire_42, N43, keyinput74);
  xor  KeyGate43 (newWire_43, N99, keyinput75);
  xnor KeyGate44 (newWire_44, N34, keyinput76);
  xor  KeyGate45 (keyNTin_Wire_1[24], N112, keyinput77);
  xor keyNTinGate_1_24(KeyNOTWire_1[12], keyinput128, keyNTin_Wire_1[24]);
  not KeyNOTGate_1_12(newWire_45, KeyNOTWire_1[12]);
  xnor KeyGate46 (keyNTin_Wire_1[25], N30, keyinput78);
  xnor keyNTinGate_1_25(KeyNOTWire_1[13], keyinput129, keyNTin_Wire_1[25]);
  not KeyNOTGate_1_13(newWire_46, KeyNOTWire_1[13]);
  xnor KeyGate47 (keyNTin_Wire_1[26], N21, keyinput79);
  xnor keyNTinGate_1_26(KeyNOTWire_1[14], keyinput130, keyNTin_Wire_1[26]);
  not KeyNOTGate_1_14(newWire_47, KeyNOTWire_1[14]);
  xnor KeyGate48 (newWire_48, N8, keyinput80);
  xor  KeyGate49 (newWire_49, N24, keyinput81);
  xor  KeyGate50 (newWire_50, N17, keyinput82);
  xnor KeyGate51 (keyNTin_Wire_1[27], N102, keyinput83);
  xnor keyNTinGate_1_27(newWire_51, keyinput131, keyNTin_Wire_1[27]);
  xor  KeyGate52 (newWire_52, N47, keyinput84);
  xor  KeyGate53 (keyNTin_Wire_1[28], N56, keyinput85);
  xnor keyNTinGate_1_28(KeyNOTWire_1[15], keyinput132, keyNTin_Wire_1[28]);
  not KeyNOTGate_1_15(newWire_53, KeyNOTWire_1[15]);
  xor  KeyGate54 (newWire_54, N79, keyinput86);
  xnor KeyGate55 (keyNTin_Wire_1[29], N40, keyinput87);
  xor keyNTinGate_1_29(KeyNOTWire_1[16], keyinput133, keyNTin_Wire_1[29]);
  not KeyNOTGate_1_16(newWire_55, KeyNOTWire_1[16]);
  xnor KeyGate56 (newWire_56, N73, keyinput88);
  xor  KeyGate57 (newWire_57, N89, keyinput89);
  xor  KeyGate58 (newWire_58, N95, keyinput90);
  xor  KeyGate59 (newWire_59, N11, keyinput91);
  xnor KeyGate60 (newWire_60, N27, keyinput92);
  xnor KeyGate61 (newWire_61, N115, keyinput93);
  xnor KeyGate62 (keyNTin_Wire_1[30], N66, keyinput94);
  xor keyNTinGate_1_30(newWire_62, keyinput134, keyNTin_Wire_1[30]);
  xor  KeyGate63 (newWire_63, N50, keyinput95);
  xor  KeyGate64 (keyNTin_Wire_1[31], N92, keyinput96);
  xor keyNTinGate_1_31(KeyNOTWire_1[17], keyinput135, keyNTin_Wire_1[31]);
  not KeyNOTGate_1_17(newWire_64, KeyNOTWire_1[17]);
  xnor KeyGate65 (newWire_65, N86, keyinput97);
  xor  KeyGate66 (newWire_66, N63, keyinput98);
  xor  KeyGate67 (newWire_67, N82, keyinput99);
  xnor KeyGate68 (keyNTin_Wire_1[32], N105, keyinput100);
  xnor keyNTinGate_1_32(KeyNOTWire_1[18], keyinput136, keyNTin_Wire_1[32]);
  not KeyNOTGate_1_18(newWire_68, KeyNOTWire_1[18]);
  xnor KeyGate69 (keyNTin_Wire_1[33], N76, keyinput101);
  xor keyNTinGate_1_33(newWire_69, keyinput137, keyNTin_Wire_1[33]);
  xnor KeyGate70 (keyNTin_Wire_1[34], N108, keyinput102);
  xor keyNTinGate_1_34(KeyNOTWire_1[19], keyinput138, keyNTin_Wire_1[34]);
  not KeyNOTGate_1_19(newWire_70, KeyNOTWire_1[19]);
  xor  KeyGate71 (keyNTin_Wire_1[35], N14, keyinput103);
  xnor keyNTinGate_1_35(newWire_71, keyinput139, keyNTin_Wire_1[35]);
  and some_function (newWire_72, newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35 );
  nand compl_function (newWire_73, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71);
  and finalAND (KeyWire_0_2, newWire_72, newWire_73);

endmodule /* AntiSAT */
