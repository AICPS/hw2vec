// Verilog File 
module top (Gid0,Gid1,Gid2,Gid3,Gid4,Gid5,Gid6,Gid7,Gid8,
Gid9,Gid10,Gid11,Gid12,Gid13,Gid14,Gid15,Gid16,Gid17,Gid18,
Gid19,Gid20,Gid21,Gid22,Gid23,Gid24,Gid25,Gid26,Gid27,Gid28,
Gid29,Gid30,Gid31,Gic0,Gic1,Gic2,Gic3,Gic4,Gic5,Gic6,
Gic7,Gr,God0,God1,God2,God3,God4,God5,God6,God7,
God8,God9,God10,God11,God12,God13,God14,God15,God16,God17,
God18,God19,God20,God21,God22,God23,God24,God25,God26,God27,
God28,God29,God30,God31,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,
keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,
keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,
keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,keyinput35,
keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,keyinput45,
keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,keyinput55,
keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,keyinput65,
keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,keyinput75,
keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,keyinput85,
keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,keyinput95,
keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,keyinput105,
keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,keyinput115,
keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,keyinput125,
keyinput126,keyinput127,keyinput128,keyinput129,keyinput130,keyinput131,keyinput132,keyinput133,keyinput134,keyinput135,
keyinput136,keyinput137,keyinput138,keyinput139,keyinput140,keyinput141,keyinput142,keyinput143,keyinput144,keyinput145,
keyinput146,keyinput147,keyinput148,keyinput149,keyinput150,keyinput151,keyinput152,keyinput153,keyinput154,keyinput155,
keyinput156,keyinput157,keyinput158,keyinput159,keyinput160,keyinput161,keyinput162,keyinput163,keyinput164,keyinput165,
keyinput166,keyinput167,keyinput168,keyinput169,keyinput170,keyinput171,keyinput172,keyinput173,keyinput174,keyinput175,
keyinput176,keyinput177,keyinput178,keyinput179,keyinput180,keyinput181,keyinput182,keyinput183,keyinput184,keyinput185,
keyinput186,keyinput187,keyinput188,keyinput189,keyinput190,keyinput191,keyinput192,keyinput193,keyinput194,keyinput195,
keyinput196,keyinput197,keyinput198,keyinput199,keyinput200,keyinput201,keyinput202,keyinput203,keyinput204,keyinput205);

input Gid0,Gid1,Gid2,Gid3,Gid4,Gid5,Gid6,Gid7,Gid8,
Gid9,Gid10,Gid11,Gid12,Gid13,Gid14,Gid15,Gid16,Gid17,Gid18,
Gid19,Gid20,Gid21,Gid22,Gid23,Gid24,Gid25,Gid26,Gid27,Gid28,
Gid29,Gid30,Gid31,Gic0,Gic1,Gic2,Gic3,Gic4,Gic5,Gic6,
Gic7,Gr,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,
keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,
keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,
keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,
keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,
keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,keyinput55,keyinput56,keyinput57,
keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,keyinput65,keyinput66,keyinput67,
keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,keyinput75,keyinput76,keyinput77,
keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,keyinput85,keyinput86,keyinput87,
keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,keyinput95,keyinput96,keyinput97,
keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,keyinput105,keyinput106,keyinput107,
keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,keyinput115,keyinput116,keyinput117,
keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,keyinput125,keyinput126,keyinput127,
keyinput128,keyinput129,keyinput130,keyinput131,keyinput132,keyinput133,keyinput134,keyinput135,keyinput136,keyinput137,
keyinput138,keyinput139,keyinput140,keyinput141,keyinput142,keyinput143,keyinput144,keyinput145,keyinput146,keyinput147,
keyinput148,keyinput149,keyinput150,keyinput151,keyinput152,keyinput153,keyinput154,keyinput155,keyinput156,keyinput157,
keyinput158,keyinput159,keyinput160,keyinput161,keyinput162,keyinput163,keyinput164,keyinput165,keyinput166,keyinput167,
keyinput168,keyinput169,keyinput170,keyinput171,keyinput172,keyinput173,keyinput174,keyinput175,keyinput176,keyinput177,
keyinput178,keyinput179,keyinput180,keyinput181,keyinput182,keyinput183,keyinput184,keyinput185,keyinput186,keyinput187,
keyinput188,keyinput189,keyinput190,keyinput191,keyinput192,keyinput193,keyinput194,keyinput195,keyinput196,keyinput197,
keyinput198,keyinput199,keyinput200,keyinput201,keyinput202,keyinput203,keyinput204,keyinput205;

output God0,God1,God2,God3,God4,God5,God6,God7,God8,
God9,God10,God11,God12,God13,God14,God15,God16,God17,God18,
God19,God20,God21,God22,God23,God24,God25,God26,God27,God28,
God29,God30,God31;

wire Gxa0,Gxa1,Gxa2,Gxa3,Gxa4,Gxa5,Gxa6,Gxa7,Gxa8,
Gxa9,Gxa10,Gxa11,Gxa12,Gxa13,Gxa14,Gxa15,Gh0,Gh1,Gh2,
Gh3,Gh4,Gh5,Gh6,Gh7,Gxb0,Gxc0,Gxb1,Gxc1,Gxb2,
Gxc2,Gxb3,Gxc3,Gxb4,Gxc4,Gxb5,Gxc5,Gxb6,Gxc6,Gxb7,
Gxc7,Gf0,Gf1,Gf2,Gf3,Gf4,Gf5,Gf6,Gf7,Gxe0,
Gxe1,Gxe2,Gxe3,Gxe4,Gxe5,Gxe6,Gxe7,Gg0,Gg1,Gg2,
Gg3,Gg4,Gg5,Gg6,Gg7,Gxd0,Gxd1,Gxd2,Gxd3,Gxd4,
Gxd5,Gxd6,Gxd7,Gs0,Gs1,Gs2,Gs3,Gs4,Gs5,Gs6,
Gs7,Gy0a,Gy1a,Gy2a,Gy0b,Gy1b,Gy3b,Gy0c,Gy2c,Gy3c,
Gy1d,Gy2d,Gy3d,Gy5i,Gy7i,Gy5j,Gy6j,Gy4k,Gy7k,Gy4l,
Gy6l,Gy4a,Gy5a,Gy6a,Gy4b,Gy5b,Gy7b,Gy4c,Gy6c,Gy7c,
Gy5d,Gy6d,Gy7d,Gy1i,Gy3i,Gy1j,Gy2j,Gy0k,Gy3k,Gy0l,
Gy2l,Gt0,Gt1,Gt2,Gt3,Gt4,Gt5,Gt6,Gt7,Gu0,
Gu1,Gwa,Gwb,Gwc,Gwd,Gwe,Gwf,Gwg,Gwh,Ge0,
Ge1,Ge2,Ge3,Ge4,Ge5,Ge6,Ge7,Ge8,Ge9,Ge10,
Ge11,Ge12,Ge13,Ge14,Ge15,Ge16,Ge17,Ge18,Ge19,Ge20,
Ge21,Ge22,Ge23,Ge24,Ge25,Ge26,Ge27,Ge28,Ge29,Ge30,
Ge31,muxed0,muxed1,muxed2,muxed3,muxed4,muxed5,muxed6,muxed7,muxed8,
muxed9,muxed10,muxed11,muxed12,muxed13,muxed14,muxed15,muxed16,muxed17,muxed18,
muxed19,muxed20,muxed21,muxed22,muxed23,muxed24,muxed25,muxed26,muxed27,muxed28,
muxed29,muxed30,muxed31,muxed32,muxed33,muxed34,muxed35,muxed36,muxed37,muxed38,
muxed39,muxed40,muxed41,muxed42,muxed43,muxed44,muxed45,muxed46,muxed47,muxed48,
muxed49,muxed50,muxed51,muxed52,muxed53,muxed54,muxed55,muxed56,muxed57,muxed58,
muxed59,muxed60,muxed61,muxed62,muxed63,muxed64,muxed65,muxed66,muxed67,muxed68,
muxed69,muxed70,muxed71,muxed72,muxed73,muxed74,muxed75,muxed76,muxed77,muxed78,
muxed79,muxed80,muxed81,muxed82,muxed83,muxed84,muxed85,muxed86,muxed87,muxed88,
muxed89,muxed90,muxed91,muxed92,muxed93,muxed94,muxed95,muxed96,muxed97,muxed98,
muxed99,muxed100,muxed101,muxed102,muxed103,muxed104,muxed105,muxed106,muxed107,muxed108,
muxed109,muxed110,muxed111,muxed112,muxed113,muxed114,muxed115,muxed116,muxed117,muxed118,
muxed119,muxed120,muxed121,muxed122,muxed123,muxed124,muxed125,muxed126,muxed127,muxed128,
muxed129,muxed130,muxed131,muxed132,muxed133,muxed134,muxed135,muxed136,muxed137,muxed138,
muxed139,muxed140,muxed141,muxed142,muxed143,muxed144,muxed145,muxed146,muxed147,muxed148,
muxed149,muxed150,muxed151,muxed152,muxed153,muxed154,muxed155,muxed156,muxed157,muxed158,
muxed159,muxed160,muxed161,muxed162,muxed163,muxed164,muxed165,muxed166,muxed167,muxed168,
muxed169,muxed170,muxed171,muxed172,muxed173,muxed174,muxed175,muxed176,muxed177,muxed178,
muxed179,muxed180,muxed181,muxed182,muxed183,muxed184,muxed185,muxed186,muxed187,muxed188,
muxed189,muxed190,muxed191,muxed192,muxed193,muxed194,muxed195,muxed196,muxed197,muxed198,
muxed199,muxed200,muxed201,muxed202,muxed203,muxed204,muxed205;
xor gate_0(Gxa0,Gid0,muxed29);
xor gate_1(Gxa1,Gid2,Gid3);
xor gate_2(Gxa2,Gid4,Gid5);
xor gate_3(Gxa3,Gid6,Gid7);
xor gate_4(Gxa4,Gid8,Gid9);
xor gate_5(Gxa5,Gid10,muxed191);
xor gate_6(Gxa6,Gid12,Gid13);
xor gate_7(Gxa7,Gid14,Gid15);
xor gate_8(Gxa8,Gid16,muxed180);
xor gate_9(Gxa9,Gid18,Gid19);
xor gate_10(Gxa10,Gid20,Gid21);
xor gate_11(Gxa11,Gid22,Gid23);
xor gate_12(Gxa12,Gid24,Gid25);
xor gate_13(Gxa13,muxed77,Gid27);
xor gate_14(Gxa14,Gid28,Gid29);
xor gate_15(Gxa15,muxed154,Gid31);
and gate_16(Gh0,Gic0,Gr);
and gate_17(Gh1,Gic1,Gr);
and gate_18(Gh2,Gic2,Gr);
and gate_19(Gh3,Gic3,Gr);
and gate_20(Gh4,Gic4,Gr);
and gate_21(Gh5,Gic5,Gr);
and gate_22(Gh6,Gic6,Gr);
and gate_23(Gh7,Gic7,Gr);
xor gate_24(Gxb0,Gid0,Gid4);
xor gate_25(Gxc0,Gid8,Gid12);
xor gate_26(Gxb1,muxed29,Gid5);
xor gate_27(Gxc1,Gid9,Gid13);
xor gate_28(Gxb2,Gid2,Gid6);
xor gate_29(Gxc2,Gid10,Gid14);
xor gate_30(Gxb3,Gid3,Gid7);
xor gate_31(Gxc3,muxed191,Gid15);
xor gate_32(Gxb4,Gid16,Gid20);
xor gate_33(Gxc4,Gid24,Gid28);
xor gate_34(Gxb5,muxed180,Gid21);
xor gate_35(Gxc5,Gid25,Gid29);
xor gate_36(Gxb6,Gid18,Gid22);
xor gate_37(Gxc6,muxed77,muxed154);
xor gate_38(Gxb7,Gid19,Gid23);
xor gate_39(Gxc7,Gid27,Gid31);
xor gate_40(Gf0,Gxa0,muxed81);
xor gate_41(Gf1,Gxa2,Gxa3);
xor gate_42(Gf2,muxed65,Gxa5);
xor gate_43(Gf3,muxed40,muxed35);
xor gate_44(Gf4,muxed31,Gxa9);
xor gate_45(Gf5,Gxa10,muxed177);
xor gate_46(Gf6,muxed203,muxed159);
xor gate_47(Gf7,Gxa14,muxed205);
xor gate_48(Gxe0,Gxb0,Gxc0);
xor gate_49(Gxe1,muxed12,muxed153);
xor gate_50(Gxe2,Gxb2,Gxc2);
xor gate_51(Gxe3,Gxb3,muxed200);
xor gate_52(Gxe4,Gxb4,Gxc4);
xor gate_53(Gxe5,muxed175,Gxc5);
xor gate_54(Gxe6,Gxb6,Gxc6);
xor gate_55(Gxe7,Gxb7,Gxc7);
xor gate_56(Gg0,Gf0,Gf1);
xor gate_57(Gg1,muxed76,muxed144);
xor gate_58(Gg2,Gf0,muxed76);
xor gate_59(Gg3,Gf1,muxed144);
xor gate_60(Gg4,muxed16,muxed189);
xor gate_61(Gg5,muxed156,muxed162);
xor gate_62(Gg6,muxed16,muxed156);
xor gate_63(Gg7,muxed189,muxed162);
xor gate_64(Gxd0,muxed110,Gg4);
xor gate_65(Gxd1,muxed123,Gg5);
xor gate_66(Gxd2,Gh2,Gg6);
xor gate_67(Gxd3,Gh3,muxed186);
xor gate_68(Gxd4,Gh4,Gg0);
xor gate_69(Gxd5,Gh5,Gg1);
xor gate_70(Gxd6,muxed160,muxed74);
xor gate_71(Gxd7,muxed13,muxed47);
xor gate_72(Gs0,Gxe0,Gxd0);
xor gate_73(Gs1,muxed14,muxed143);
xor gate_74(Gs2,muxed167,Gxd2);
xor gate_75(Gs3,muxed198,muxed170);
xor gate_76(Gs4,muxed26,Gxd4);
xor gate_77(Gs5,Gxe5,Gxd5);
xor gate_78(Gs6,Gxe6,muxed72);
xor gate_79(Gs7,Gxe7,muxed45);
not gate_80(Gy0a,Gs0);
not gate_81(Gy1a,muxed140);
not gate_82(Gy2a,muxed141);
not gate_83(Gy0b,Gs0);
not gate_84(Gy1b,muxed140);
not gate_85(Gy3b,muxed195);
not gate_86(Gy0c,Gs0);
not gate_87(Gy2c,muxed141);
not gate_88(Gy3c,muxed195);
not gate_89(Gy1d,muxed140);
not gate_90(Gy2d,muxed141);
not gate_91(Gy3d,muxed195);
not gate_92(Gy5i,Gs5);
not gate_93(Gy7i,muxed44);
not gate_94(Gy5j,Gs5);
not gate_95(Gy6j,muxed85);
not gate_96(Gy4k,Gs4);
not gate_97(Gy7k,muxed44);
not gate_98(Gy4l,Gs4);
not gate_99(Gy6l,muxed85);
not gate_100(Gy4a,Gs4);
not gate_101(Gy5a,Gs5);
not gate_102(Gy6a,muxed85);
not gate_103(Gy4b,Gs4);
not gate_104(Gy5b,Gs5);
not gate_105(Gy7b,muxed44);
not gate_106(Gy4c,Gs4);
not gate_107(Gy6c,muxed85);
not gate_108(Gy7c,muxed44);
not gate_109(Gy5d,Gs5);
not gate_110(Gy6d,muxed85);
not gate_111(Gy7d,muxed44);
not gate_112(Gy1i,muxed140);
not gate_113(Gy3i,muxed195);
not gate_114(Gy1j,muxed140);
not gate_115(Gy2j,muxed141);
not gate_116(Gy0k,Gs0);
not gate_117(Gy3k,muxed195);
not gate_118(Gy0l,Gs0);
not gate_119(Gy2l,muxed141);
and gate_120(Gt0,Gy0a,muxed152,muxed126,muxed195);
and gate_121(Gt1,muxed184,Gy1b,muxed141,Gy3b);
and gate_122(Gt2,muxed136,muxed140,Gy2c,Gy3c);
and gate_123(Gt3,Gs0,muxed84,Gy2d,Gy3d);
and gate_124(Gt4,Gy4a,Gy5a,muxed62,muxed44);
and gate_125(Gt5,muxed101,Gy5b,muxed85,Gy7b);
and gate_126(Gt6,Gy4c,Gs5,Gy6c,muxed11);
and gate_127(Gt7,Gs4,Gy5d,Gy6d,Gy7d);
or gate_128(Gu0,muxed182,muxed19,muxed7,Gt3);
or gate_129(Gu1,muxed92,muxed111,muxed164,Gt7);
and gate_130(Gwa,Gs4,muxed129,muxed85,muxed199,muxed119);
and gate_131(Gwb,Gs4,Gy5j,muxed146,muxed44,muxed119);
and gate_132(Gwc,Gy4k,Gs5,muxed85,Gy7k,muxed119);
and gate_133(Gwd,muxed89,Gs5,Gy6l,muxed44,muxed119);
and gate_134(Gwe,Gs0,Gy1i,muxed141,Gy3i,muxed108);
and gate_135(Gwf,Gs0,muxed114,Gy2j,muxed195,muxed108);
and gate_136(Gwg,muxed105,muxed140,muxed141,Gy3k,muxed108);
and gate_137(Gwh,Gy0l,muxed140,Gy2l,muxed195,muxed108);
and gate_138(Ge0,Gs0,muxed51);
and gate_139(Ge1,muxed140,muxed51);
and gate_140(Ge2,muxed141,muxed51);
and gate_141(Ge3,muxed195,muxed51);
and gate_142(Ge4,Gs0,Gwb);
and gate_143(Ge5,muxed140,Gwb);
and gate_144(Ge6,muxed141,Gwb);
and gate_145(Ge7,muxed195,Gwb);
and gate_146(Ge8,Gs0,Gwc);
and gate_147(Ge9,muxed140,Gwc);
and gate_148(Ge10,muxed141,Gwc);
and gate_149(Ge11,muxed195,Gwc);
and gate_150(Ge12,Gs0,muxed98);
and gate_151(Ge13,muxed140,muxed98);
and gate_152(Ge14,muxed141,muxed98);
and gate_153(Ge15,muxed195,muxed98);
and gate_154(Ge16,Gs4,Gwe);
and gate_155(Ge17,Gs5,Gwe);
and gate_156(Ge18,muxed85,Gwe);
and gate_157(Ge19,muxed44,Gwe);
and gate_158(Ge20,Gs4,muxed54);
and gate_159(Ge21,Gs5,muxed54);
and gate_160(Ge22,muxed85,muxed54);
and gate_161(Ge23,muxed44,muxed54);
and gate_162(Ge24,Gs4,muxed36);
and gate_163(Ge25,Gs5,muxed36);
and gate_164(Ge26,muxed85,muxed36);
and gate_165(Ge27,muxed44,muxed36);
and gate_166(Ge28,Gs4,muxed106);
and gate_167(Ge29,Gs5,muxed106);
and gate_168(Ge30,muxed85,muxed106);
and gate_169(Ge31,muxed44,muxed106);
xor gate_170(God0,Gid0,muxed75);
xor gate_171(God1,muxed29,muxed201);
xor gate_172(God2,Gid2,Ge2);
xor gate_173(God3,Gid3,Ge3);
xor gate_174(God4,Gid4,Ge4);
xor gate_175(God5,Gid5,Ge5);
xor gate_176(God6,Gid6,Ge6);
xor gate_177(God7,Gid7,Ge7);
xor gate_178(God8,Gid8,Ge8);
xor gate_179(God9,Gid9,muxed55);
xor gate_180(God10,Gid10,Ge10);
xor gate_181(God11,muxed191,Ge11);
xor gate_182(God12,Gid12,Ge12);
xor gate_183(God13,Gid13,muxed127);
xor gate_184(God14,Gid14,muxed96);
xor gate_185(God15,Gid15,muxed21);
xor gate_186(God16,Gid16,Ge16);
xor gate_187(God17,muxed180,Ge17);
xor gate_188(God18,Gid18,muxed82);
xor gate_189(God19,Gid19,Ge19);
xor gate_190(God20,Gid20,Ge20);
xor gate_191(God21,Gid21,Ge21);
xor gate_192(God22,Gid22,Ge22);
xor gate_193(God23,Gid23,muxed183);
xor gate_194(God24,Gid24,Ge24);
xor gate_195(God25,Gid25,Ge25);
xor gate_196(God26,muxed77,Ge26);
xor gate_197(God27,Gid27,muxed197);
xor gate_198(God28,Gid28,Ge28);
xor gate_199(God29,Gid29,muxed71);
xor gate_200(God30,muxed154,Ge30);
xor gate_201(God31,Gid31,muxed150);
assign muxed0 = keyinput0 ? Gid1 : muxed161;
assign muxed1 = keyinput1 ? muxed57 : Ge16;
assign muxed2 = keyinput2 ? Ge9 : muxed57;
assign muxed3 = keyinput3 ? muxed97 : muxed127;
assign muxed4 = keyinput4 ? muxed50 : muxed97;
assign muxed5 = keyinput5 ? muxed99 : Gy6c;
assign muxed6 = keyinput6 ? muxed120 : muxed11;
assign muxed7 = keyinput7 ? muxed139 : Ge24;
assign muxed8 = keyinput8 ? muxed38 : muxed139;
assign muxed9 = keyinput9 ? muxed25 : Gf1;
assign muxed10 = keyinput10 ? Gxe1 : Gxb0;
assign muxed11 = keyinput11 ? Gy7c : Gxe1;
assign muxed12 = keyinput12 ? Gxb1 : Gt3;
assign muxed13 = keyinput13 ? Gh7 : Gxb1;
assign muxed14 = keyinput14 ? muxed171 : muxed15;
assign muxed15 = keyinput15 ? muxed131 : Gy7b;
assign muxed16 = keyinput16 ? Gf4 : muxed131;
assign muxed17 = keyinput17 ? muxed30 : Gxe0;
assign muxed18 = keyinput18 ? muxed1 : muxed36;
assign muxed19 = keyinput19 ? Gt1 : muxed1;
assign muxed20 = keyinput20 ? God15 : muxed71;
assign muxed21 = keyinput21 ? muxed79 : muxed171;
assign muxed22 = keyinput22 ? muxed32 : muxed79;
assign muxed23 = keyinput23 ? Ge13 : muxed44;
assign muxed24 = keyinput24 ? muxed9 : muxed54;
assign muxed25 = keyinput25 ? muxed90 : Gy1b;
assign muxed26 = keyinput26 ? Gxe4 : muxed90;
assign muxed27 = keyinput27 ? Gxe2 : muxed131;
assign muxed28 = keyinput28 ? God1 : Gy2c;
assign muxed29 = keyinput29 ? muxed17 : Gxa14;
assign muxed30 = keyinput30 ? muxed41 : Ge2;
assign muxed31 = keyinput31 ? Gxa8 : muxed41;
assign muxed32 = keyinput32 ? muxed0 : muxed146;
assign muxed33 = keyinput33 ? muxed113 : muxed0;
assign muxed34 = keyinput34 ? muxed18 : muxed162;
assign muxed35 = keyinput35 ? muxed64 : muxed18;
assign muxed36 = keyinput36 ? Gwg : Gy2j;
assign muxed37 = keyinput37 ? muxed137 : muxed153;
assign muxed38 = keyinput38 ? muxed179 : muxed54;
assign muxed39 = keyinput39 ? Gxa11 : muxed179;
assign muxed40 = keyinput40 ? Gxa6 : muxed41;
assign muxed41 = keyinput41 ? muxed66 : muxed32;
assign muxed42 = keyinput42 ? muxed3 : muxed82;
assign muxed43 = keyinput43 ? muxed23 : Ge13;
assign muxed44 = keyinput44 ? Gs7 : muxed167;
assign muxed45 = keyinput45 ? Gxd7 : muxed141;
assign muxed46 = keyinput46 ? muxed204 : Gxd7;
assign muxed47 = keyinput47 ? muxed93 : muxed51;
assign muxed48 = keyinput48 ? Gxd1 : muxed93;
assign muxed49 = keyinput49 ? muxed149 : Gf0;
assign muxed50 = keyinput50 ? Gf3 : Gy3b;
assign muxed51 = keyinput51 ? Gwa : Gf3;
assign muxed52 = keyinput52 ? muxed70 : muxed53;
assign muxed53 = keyinput53 ? God9 : Gy5d;
assign muxed54 = keyinput54 ? Gwf : God9;
assign muxed55 = keyinput55 ? muxed73 : Gwf;
assign muxed56 = keyinput56 ? Gh0 : muxed73;
assign muxed57 = keyinput57 ? muxed20 : Gf4;
assign muxed58 = keyinput58 ? Ge29 : Gxb0;
assign muxed59 = keyinput59 ? muxed133 : Ge12;
assign muxed60 = keyinput60 ? muxed109 : muxed45;
assign muxed61 = keyinput61 ? Gt4 : muxed133;
assign muxed62 = keyinput62 ? muxed63 : Gt4;
assign muxed63 = keyinput63 ? Gy6a : muxed146;
assign muxed64 = keyinput64 ? Gxa7 : Gy6a;
assign muxed65 = keyinput65 ? Gxa4 : muxed66;
assign muxed66 = keyinput66 ? muxed78 : Ge19;
assign muxed67 = keyinput67 ? muxed80 : Gxe1;
assign muxed68 = keyinput68 ? muxed83 : Gy2c;
assign muxed69 = keyinput69 ? muxed158 : muxed156;
assign muxed70 = keyinput70 ? Gs6 : Gxe4;
assign muxed71 = keyinput71 ? muxed58 : Gs6;
assign muxed72 = keyinput72 ? muxed166 : Gy6a;
assign muxed73 = keyinput73 ? muxed2 : muxed166;
assign muxed74 = keyinput74 ? Gg2 : muxed0;
assign muxed75 = keyinput75 ? Ge0 : Gg2;
assign muxed76 = keyinput76 ? Gf2 : Gy6a;
assign muxed77 = keyinput77 ? Gid26 : muxed78;
assign muxed78 = keyinput78 ? muxed22 : muxed53;
assign muxed79 = keyinput79 ? muxed67 : Gxb3;
assign muxed80 = keyinput80 ? muxed42 : Gs0;
assign muxed81 = keyinput81 ? Gxa1 : muxed42;
assign muxed82 = keyinput82 ? muxed68 : Gy3d;
assign muxed83 = keyinput83 ? Ge18 : Gg5;
assign muxed84 = keyinput84 ? Gy1d : Ge18;
assign muxed85 = keyinput85 ? muxed155 : muxed110;
assign muxed86 = keyinput86 ? muxed157 : Gy2c;
assign muxed87 = keyinput87 ? Gxa13 : muxed161;
assign muxed88 = keyinput88 ? muxed202 : Gxa13;
assign muxed89 = keyinput89 ? Gy4l : muxed90;
assign muxed90 = keyinput90 ? Gs1 : muxed45;
assign muxed91 = keyinput91 ? muxed48 : Gy3i;
assign muxed92 = keyinput92 ? muxed61 : muxed48;
assign muxed93 = keyinput93 ? Gg3 : muxed54;
assign muxed94 = keyinput94 ? muxed147 : muxed129;
assign muxed95 = keyinput95 ? muxed4 : Ge7;
assign muxed96 = keyinput96 ? Ge14 : muxed4;
assign muxed97 = keyinput97 ? muxed192 : muxed199;
assign muxed98 = keyinput98 ? muxed5 : muxed201;
assign muxed99 = keyinput99 ? muxed132 : muxed127;
assign muxed100 = keyinput100 ? Gy5i : muxed132;
assign muxed101 = keyinput101 ? muxed178 : muxed102;
assign muxed102 = keyinput102 ? God31 : muxed184;
assign muxed103 = keyinput103 ? muxed122 : God31;
assign muxed104 = keyinput104 ? Ge31 : muxed20;
assign muxed105 = keyinput105 ? Gy0k : Ge31;
assign muxed106 = keyinput106 ? muxed59 : muxed5;
assign muxed107 = keyinput107 ? Gwh : muxed141;
assign muxed108 = keyinput108 ? muxed60 : Gxb6;
assign muxed109 = keyinput109 ? Gu1 : Ge6;
assign muxed110 = keyinput110 ? muxed56 : Gu1;
assign muxed111 = keyinput111 ? muxed33 : Gwg;
assign muxed112 = keyinput112 ? muxed172 : muxed33;
assign muxed113 = keyinput113 ? Gt5 : Gy2j;
assign muxed114 = keyinput114 ? Gy1j : Gt5;
assign muxed115 = keyinput115 ? muxed135 : muxed144;
assign muxed116 = keyinput116 ? muxed145 : Ge0;
assign muxed117 = keyinput117 ? muxed130 : Ge12;
assign muxed118 = keyinput118 ? Gwd : muxed133;
assign muxed119 = keyinput119 ? muxed6 : Gy0l;
assign muxed120 = keyinput120 ? muxed103 : muxed67;
assign muxed121 = keyinput121 ? Gy0c : muxed103;
assign muxed122 = keyinput122 ? muxed181 : Gg6;
assign muxed123 = keyinput123 ? Gh1 : muxed181;
assign muxed124 = keyinput124 ? muxed151 : muxed184;
assign muxed125 = keyinput125 ? muxed95 : muxed151;
assign muxed126 = keyinput126 ? Gy2a : Gs6;
assign muxed127 = keyinput127 ? muxed43 : Gy2a;
assign muxed128 = keyinput128 ? muxed121 : muxed129;
assign muxed129 = keyinput129 ? muxed117 : Ge25;
assign muxed130 = keyinput130 ? muxed100 : muxed102;
assign muxed131 = keyinput131 ? muxed28 : muxed100;
assign muxed132 = keyinput132 ? muxed118 : muxed43;
assign muxed133 = keyinput133 ? muxed107 : Gxd4;
assign muxed134 = keyinput134 ? muxed142 : muxed58;
assign muxed135 = keyinput135 ? muxed37 : muxed80;
assign muxed136 = keyinput136 ? muxed128 : muxed37;
assign muxed137 = keyinput137 ? muxed8 : muxed139;
assign muxed138 = keyinput138 ? muxed163 : muxed8;
assign muxed139 = keyinput139 ? Gt2 : muxed108;
assign muxed140 = keyinput140 ? muxed24 : muxed141;
assign muxed141 = keyinput141 ? muxed134 : Ge7;
assign muxed142 = keyinput142 ? muxed115 : muxed81;
assign muxed143 = keyinput143 ? muxed91 : muxed115;
assign muxed144 = keyinput144 ? muxed116 : Gxa13;
assign muxed145 = keyinput145 ? muxed94 : muxed26;
assign muxed146 = keyinput146 ? Gy6j : muxed94;
assign muxed147 = keyinput147 ? muxed49 : Gy3i;
assign muxed148 = keyinput148 ? Gy0b : muxed49;
assign muxed149 = keyinput149 ? muxed125 : Gy2d;
assign muxed150 = keyinput150 ? muxed104 : muxed125;
assign muxed151 = keyinput151 ? Gt0 : Gxa9;
assign muxed152 = keyinput152 ? Gy1a : muxed104;
assign muxed153 = keyinput153 ? muxed187 : Gy1a;
assign muxed154 = keyinput154 ? Gid30 : muxed155;
assign muxed155 = keyinput155 ? muxed69 : Gf4;
assign muxed156 = keyinput156 ? muxed86 : Gwg;
assign muxed157 = keyinput157 ? Gf6 : Gg2;
assign muxed158 = keyinput158 ? muxed52 : Gf6;
assign muxed159 = keyinput159 ? muxed87 : Gxb3;
assign muxed160 = keyinput160 ? Gh6 : muxed87;
assign muxed161 = keyinput161 ? muxed34 : Gxb2;
assign muxed162 = keyinput162 ? muxed138 : Gy6l;
assign muxed163 = keyinput163 ? Gf7 : Gf1;
assign muxed164 = keyinput164 ? Gt6 : Gf7;
assign muxed165 = keyinput165 ? Gxa15 : muxed154;
assign muxed166 = keyinput166 ? Gxd6 : Gxa15;
assign muxed167 = keyinput167 ? muxed27 : muxed192;
assign muxed168 = keyinput168 ? muxed193 : Gxa10;
assign muxed169 = keyinput169 ? muxed196 : muxed6;
assign muxed170 = keyinput170 ? muxed112 : muxed199;
assign muxed171 = keyinput171 ? muxed10 : muxed112;
assign muxed172 = keyinput172 ? muxed185 : muxed10;
assign muxed173 = keyinput173 ? muxed148 : muxed185;
assign muxed174 = keyinput174 ? muxed188 : Gxc5;
assign muxed175 = keyinput175 ? muxed190 : muxed188;
assign muxed176 = keyinput176 ? muxed194 : muxed190;
assign muxed177 = keyinput177 ? muxed39 : muxed9;
assign muxed178 = keyinput178 ? Gy4b : muxed39;
assign muxed179 = keyinput179 ? Gs2 : Gs1;
assign muxed180 = keyinput180 ? Gid17 : muxed181;
assign muxed181 = keyinput181 ? Gu0 : Gy2c;
assign muxed182 = keyinput182 ? muxed124 : Gh4;
assign muxed183 = keyinput183 ? Ge23 : muxed124;
assign muxed184 = keyinput184 ? muxed173 : Gy0b;
assign muxed185 = keyinput185 ? Gxd3 : Gxb6;
assign muxed186 = keyinput186 ? muxed174 : Ge26;
assign muxed187 = keyinput187 ? Gxc1 : muxed174;
assign muxed188 = keyinput188 ? Gg7 : Ge4;
assign muxed189 = keyinput189 ? muxed176 : muxed86;
assign muxed190 = keyinput190 ? Gxb5 : Gg2;
assign muxed191 = keyinput191 ? Gid11 : muxed192;
assign muxed192 = keyinput192 ? muxed168 : Gt0;
assign muxed193 = keyinput193 ? Ge15 : muxed132;
assign muxed194 = keyinput194 ? Gf5 : Ge15;
assign muxed195 = keyinput195 ? muxed169 : Gy2c;
assign muxed196 = keyinput196 ? Gs3 : Gxa1;
assign muxed197 = keyinput197 ? Ge27 : Gs3;
assign muxed198 = keyinput198 ? Gxe3 : muxed178;
assign muxed199 = keyinput199 ? Gy7i : Gxe3;
assign muxed200 = keyinput200 ? muxed88 : muxed123;
assign muxed201 = keyinput201 ? Ge1 : muxed88;
assign muxed202 = keyinput202 ? muxed46 : muxed70;
assign muxed203 = keyinput203 ? Gxa12 : muxed46;
assign muxed204 = keyinput204 ? Gxc3 : Gxe5;
assign muxed205 = keyinput205 ? muxed165 : Gxc3;
endmodule
