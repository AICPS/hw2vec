`timescale 1ns / 1ps
// Verilog
// c432
// Ninputs 36
// Noutputs 7
// NtotalGates 160
// NOT1 40
// NAND2 64
// NOR2 19
// AND9 3
// XOR2 18
// NAND4 14
// AND8 1
// NAND3 1

module top (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
                  N430,N431,N432,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
                  keyinput60, keyinput61, keyinput62, keyinput63,
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
        keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
        keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
        keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
        keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
        keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
                  keyinput134, keyinput135,
        keyinput136, keyinput137, keyinput138, keyinput139, keyinput140,
        keyinput141, keyinput142, keyinput143, keyinput144, keyinput145,
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150,
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155,
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160,
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165,
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170,
        keyinput171);

  input keyinput136, keyinput137, keyinput138, keyinput139, keyinput140;
  input keyinput141, keyinput142, keyinput143, keyinput144, keyinput145;
  input keyinput146, keyinput147, keyinput148, keyinput149, keyinput150;
  input keyinput151, keyinput152, keyinput153, keyinput154, keyinput155;
  input keyinput156, keyinput157, keyinput158, keyinput159, keyinput160;
  input keyinput161, keyinput162, keyinput163, keyinput164, keyinput165;
  input keyinput166, keyinput167, keyinput168, keyinput169, keyinput170;
  input keyinput171;


  input keyinput64, keyinput65, keyinput66, keyinput67, keyinput68;
  input keyinput69, keyinput70, keyinput71, keyinput72, keyinput73;
  input keyinput74, keyinput75, keyinput76, keyinput77, keyinput78;
  input keyinput79, keyinput80, keyinput81, keyinput82, keyinput83;
  input keyinput84, keyinput85, keyinput86, keyinput87, keyinput88;
  input keyinput89, keyinput90, keyinput91, keyinput92, keyinput93;
  input keyinput94, keyinput95, keyinput96, keyinput97, keyinput98;
  input keyinput99, keyinput100, keyinput101, keyinput102, keyinput103;
  input keyinput104, keyinput105, keyinput106, keyinput107, keyinput108;
  input keyinput109, keyinput110, keyinput111, keyinput112, keyinput113;
  input keyinput114, keyinput115, keyinput116, keyinput117, keyinput118;
  input keyinput119, keyinput120, keyinput121, keyinput122, keyinput123;
  input keyinput124, keyinput125, keyinput126, keyinput127, keyinput128;
  input keyinput129, keyinput130, keyinput131, keyinput132, keyinput133;
  input keyinput134, keyinput135;

  wire KeyWire_0_1 , KeyWire_0_2;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31, keyinput32, keyinput33, keyinput34;
  input keyinput35, keyinput36, keyinput37, keyinput38, keyinput39;
  input keyinput40, keyinput41, keyinput42, keyinput43, keyinput44;
  input keyinput45, keyinput46, keyinput47, keyinput48, keyinput49;
  input keyinput50, keyinput51, keyinput52, keyinput53, keyinput54;
  input keyinput55, keyinput56, keyinput57, keyinput58, keyinput59;
  input keyinput60, keyinput61, keyinput62, keyinput63;

  wire [0:63] keyinput_Wire_0;
  wire [0:26] KeyNOTWire_0;

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;

output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429;

  not NOT1_1 (keyinput_Wire_0[0], N1);
  xor keyGate_0_0(KeyNOTWire_0[0], keyinput0, keyinput_Wire_0[0]);
  not KeyNOTGate_0_0(N118, KeyNOTWire_0[0]);
  not NOT1_2 (keyinput_Wire_0[1], N4);
  xnor keyGate_0_1(KeyNOTWire_0[1], keyinput1, keyinput_Wire_0[1]);
  not KeyNOTGate_0_1(N119, KeyNOTWire_0[1]);
  not NOT1_3 (keyinput_Wire_0[2], N11);
  xor keyGate_0_2(N122, keyinput2, keyinput_Wire_0[2]);
  not NOT1_4 (keyinput_Wire_0[3], N17);
  xor keyGate_0_3(KeyNOTWire_0[2], keyinput3, keyinput_Wire_0[3]);
  not KeyNOTGate_0_2(N123, KeyNOTWire_0[2]);
  not NOT1_5 (keyinput_Wire_0[4], N24);
  xor keyGate_0_4(N126, keyinput4, keyinput_Wire_0[4]);
  not NOT1_6 (keyinput_Wire_0[5], N30);
  xor keyGate_0_5(N127, keyinput5, keyinput_Wire_0[5]);
  not NOT1_7 (keyinput_Wire_0[6], N37);
  xnor keyGate_0_6(N130, keyinput6, keyinput_Wire_0[6]);
  not NOT1_8 (keyinput_Wire_0[7], N43);
  xnor keyGate_0_7(KeyNOTWire_0[3], keyinput7, keyinput_Wire_0[7]);
  not KeyNOTGate_0_3(N131, KeyNOTWire_0[3]);
  not NOT1_9 (keyinput_Wire_0[8], N50);
  xnor keyGate_0_8(KeyNOTWire_0[4], keyinput8, keyinput_Wire_0[8]);
  not KeyNOTGate_0_4(N134, KeyNOTWire_0[4]);
  not NOT1_10 (keyinput_Wire_0[9], N56);
  xnor keyGate_0_9(N135, keyinput9, keyinput_Wire_0[9]);
  not NOT1_11 (keyinput_Wire_0[10], N63);
  xnor keyGate_0_10(KeyNOTWire_0[5], keyinput10, keyinput_Wire_0[10]);
  not KeyNOTGate_0_5(N138, KeyNOTWire_0[5]);
  not NOT1_12 (keyinput_Wire_0[11], N69);
  xor keyGate_0_11(N139, keyinput11, keyinput_Wire_0[11]);
  not NOT1_13 (keyinput_Wire_0[12], N76);
  xnor keyGate_0_12(N142, keyinput12, keyinput_Wire_0[12]);
  not NOT1_14 (keyinput_Wire_0[13], N82);
  xnor keyGate_0_13(N143, keyinput13, keyinput_Wire_0[13]);
  not NOT1_15 (keyinput_Wire_0[14], N89);
  xor keyGate_0_14(KeyNOTWire_0[6], keyinput14, keyinput_Wire_0[14]);
  not KeyNOTGate_0_6(N146, KeyNOTWire_0[6]);
  not NOT1_16 (keyinput_Wire_0[15], N95);
  xnor keyGate_0_15(KeyNOTWire_0[7], keyinput15, keyinput_Wire_0[15]);
  not KeyNOTGate_0_7(N147, KeyNOTWire_0[7]);
  not NOT1_17 (keyinput_Wire_0[16], N102);
  xnor keyGate_0_16(KeyNOTWire_0[8], keyinput16, keyinput_Wire_0[16]);
  not KeyNOTGate_0_8(N150, KeyNOTWire_0[8]);
  not NOT1_18 (keyinput_Wire_0[17], N108);
  xor keyGate_0_17(N151, keyinput17, keyinput_Wire_0[17]);
  nand NAND2_19 (keyinput_Wire_0[18], N118, N4);
  xor keyGate_0_18(N154, keyinput18, keyinput_Wire_0[18]);
  nor NOR2_20 (keyinput_Wire_0[19], N8, N119);
  xnor keyGate_0_19(N157, keyinput19, keyinput_Wire_0[19]);
  nor NOR2_21 (keyinput_Wire_0[20], N14, N119);
  xor keyGate_0_20(N158, keyinput20, keyinput_Wire_0[20]);
  nand NAND2_22 (keyinput_Wire_0[21], N122, N17);
  xor keyGate_0_21(KeyNOTWire_0[9], keyinput21, keyinput_Wire_0[21]);
  not KeyNOTGate_0_9(N159, KeyNOTWire_0[9]);
  nand NAND2_23 (keyinput_Wire_0[22], N126, N30);
  xnor keyGate_0_22(N162, keyinput22, keyinput_Wire_0[22]);
  nand NAND2_24 (keyinput_Wire_0[23], N130, N43);
  xnor keyGate_0_23(N165, keyinput23, keyinput_Wire_0[23]);
  nand NAND2_25 (keyinput_Wire_0[24], N134, N56);
  xor keyGate_0_24(N168, keyinput24, keyinput_Wire_0[24]);
  nand NAND2_26 (keyinput_Wire_0[25], N138, N69);
  xnor keyGate_0_25(KeyNOTWire_0[10], keyinput25, keyinput_Wire_0[25]);
  not KeyNOTGate_0_10(N171, KeyNOTWire_0[10]);
  nand NAND2_27 (keyinput_Wire_0[26], N142, N82);
  xor keyGate_0_26(N174, keyinput26, keyinput_Wire_0[26]);
  nand NAND2_28 (keyinput_Wire_0[27], N146, N95);
  xor keyGate_0_27(N177, keyinput27, keyinput_Wire_0[27]);
  nand NAND2_29 (keyinput_Wire_0[28], N150, N108);
  xor keyGate_0_28(KeyNOTWire_0[11], keyinput28, keyinput_Wire_0[28]);
  not KeyNOTGate_0_11(N180, KeyNOTWire_0[11]);
  nor NOR2_30 (keyinput_Wire_0[29], N21, N123);
  xnor keyGate_0_29(N183, keyinput29, keyinput_Wire_0[29]);
nor NOR2_31 (N184, N27, N123);
nor NOR2_32 (N185, N34, N127);
  nor NOR2_33 (keyinput_Wire_0[30], N40, N127);
  xor keyGate_0_30(N186, keyinput30, keyinput_Wire_0[30]);
nor NOR2_34 (N187, N47, N131);
  nor NOR2_35 (keyinput_Wire_0[31], N53, N131);
  xor keyGate_0_31(KeyNOTWire_0[12], keyinput31, keyinput_Wire_0[31]);
  not KeyNOTGate_0_12(N188, KeyNOTWire_0[12]);
  nor NOR2_36 (keyinput_Wire_0[32], N60, N135);
  xnor keyGate_0_32(KeyNOTWire_0[13], keyinput32, keyinput_Wire_0[32]);
  not KeyNOTGate_0_13(N189, KeyNOTWire_0[13]);
  nor NOR2_37 (keyinput_Wire_0[33], N66, N135);
  xor keyGate_0_33(N190, keyinput33, keyinput_Wire_0[33]);
  nor NOR2_38 (keyinput_Wire_0[34], N73, N139);
  xor keyGate_0_34(N191, keyinput34, keyinput_Wire_0[34]);
nor NOR2_39 (N192, N79, N139);
  nor NOR2_40 (keyinput_Wire_0[35], N86, N143);
  xnor keyGate_0_35(N193, keyinput35, keyinput_Wire_0[35]);
nor NOR2_41 (N194, N92, N143);
  nor NOR2_42 (keyinput_Wire_0[36], N99, N147);
  xor keyGate_0_36(KeyNOTWire_0[14], keyinput36, keyinput_Wire_0[36]);
  not KeyNOTGate_0_14(N195, KeyNOTWire_0[14]);
  nor NOR2_43 (keyinput_Wire_0[37], N105, N147);
  xnor keyGate_0_37(N196, keyinput37, keyinput_Wire_0[37]);
  nor NOR2_44 (keyinput_Wire_0[38], N112, N151);
  xor keyGate_0_38(N197, keyinput38, keyinput_Wire_0[38]);
nor NOR2_45 (N198, N115, N151);
  and AND9_46 (keyinput_Wire_0[39], N154, N159, N162, N165, N168, N171, N174, N177, N180);
  xnor keyGate_0_39(N199, keyinput39, keyinput_Wire_0[39]);
  not NOT1_47 (keyinput_Wire_0[40], N199);
  xor keyGate_0_40(N203, keyinput40, keyinput_Wire_0[40]);
not NOT1_48 (N213, N199);
not NOT1_49 (N223, N199);
  xor XOR2_50 (keyinput_Wire_0[41], N203, N154);
  xor keyGate_0_41(N224, keyinput41, keyinput_Wire_0[41]);
  xor XOR2_51 (keyinput_Wire_0[42], N203, N159);
  xor keyGate_0_42(KeyNOTWire_0[15], keyinput42, keyinput_Wire_0[42]);
  not KeyNOTGate_0_15(N227, KeyNOTWire_0[15]);
  xor XOR2_52 (keyinput_Wire_0[43], N203, N162);
  xor keyGate_0_43(KeyNOTWire_0[16], keyinput43, keyinput_Wire_0[43]);
  not KeyNOTGate_0_16(N230, KeyNOTWire_0[16]);
  xor XOR2_53 (keyinput_Wire_0[44], N203, N165);
  xnor keyGate_0_44(KeyNOTWire_0[17], keyinput44, keyinput_Wire_0[44]);
  not KeyNOTGate_0_17(N233, KeyNOTWire_0[17]);
  xor XOR2_54 (keyinput_Wire_0[45], N203, N168);
  xor keyGate_0_45(KeyNOTWire_0[18], keyinput45, keyinput_Wire_0[45]);
  not KeyNOTGate_0_18(N236, KeyNOTWire_0[18]);
  xor XOR2_55 (keyinput_Wire_0[46], N203, N171);
  xnor keyGate_0_46(N239, keyinput46, keyinput_Wire_0[46]);
nand NAND2_56 (N242, N1, N213);
  xor XOR2_57 (keyinput_Wire_0[47], N203, N174);
  xnor keyGate_0_47(N243, keyinput47, keyinput_Wire_0[47]);
nand NAND2_58 (N246, N213, N11);
  xor XOR2_59 (keyinput_Wire_0[48], N203, N177);
  xor keyGate_0_48(N247, keyinput48, keyinput_Wire_0[48]);
nand NAND2_60 (N250, N213, N24);
  xor XOR2_61 (keyinput_Wire_0[49], N203, N180);
  xor keyGate_0_49(N251, keyinput49, keyinput_Wire_0[49]);
nand NAND2_62 (N254, N213, N37);
nand NAND2_63 (N255, N213, N50);
nand NAND2_64 (N256, N213, N63);
nand NAND2_65 (N257, N213, N76);
nand NAND2_66 (N258, N213, N89);
nand NAND2_67 (N259, N213, N102);
  nand NAND2_68 (keyinput_Wire_0[50], N224, N157);
  xnor keyGate_0_50(KeyNOTWire_0[19], keyinput50, keyinput_Wire_0[50]);
  not KeyNOTGate_0_19(N260, KeyNOTWire_0[19]);
nand NAND2_69 (N263, N224, N158);
nand NAND2_70 (N264, N227, N183);
  nand NAND2_71 (keyinput_Wire_0[51], N230, N185);
  xnor keyGate_0_51(KeyNOTWire_0[20], keyinput51, keyinput_Wire_0[51]);
  not KeyNOTGate_0_20(N267, KeyNOTWire_0[20]);
  nand NAND2_72 (keyinput_Wire_0[52], N233, N187);
  xnor keyGate_0_52(N270, keyinput52, keyinput_Wire_0[52]);
  nand NAND2_73 (keyinput_Wire_0[53], N236, N189);
  xnor keyGate_0_53(N273, keyinput53, keyinput_Wire_0[53]);
  nand NAND2_74 (keyinput_Wire_0[54], N239, N191);
  xor keyGate_0_54(KeyNOTWire_0[21], keyinput54, keyinput_Wire_0[54]);
  not KeyNOTGate_0_21(N276, KeyNOTWire_0[21]);
  nand NAND2_75 (keyinput_Wire_0[55], N243, N193);
  xor keyGate_0_55(KeyNOTWire_0[22], keyinput55, keyinput_Wire_0[55]);
  not KeyNOTGate_0_22(N279, KeyNOTWire_0[22]);
  nand NAND2_76 (keyinput_Wire_0[56], N247, N195);
  xnor keyGate_0_56(KeyNOTWire_0[23], keyinput56, keyinput_Wire_0[56]);
  not KeyNOTGate_0_23(N282, KeyNOTWire_0[23]);
nand NAND2_77 (N285, N251, N197);
nand NAND2_78 (N288, N227, N184);
nand NAND2_79 (N289, N230, N186);
nand NAND2_80 (N290, N233, N188);
nand NAND2_81 (N291, N236, N190);
nand NAND2_82 (N292, N239, N192);
nand NAND2_83 (N293, N243, N194);
nand NAND2_84 (N294, N247, N196);
nand NAND2_85 (N295, N251, N198);
and AND9_86 (N296, N260, N264, N267, N270, N273, N276, N279, N282, N285);
  not NOT1_87 (keyinput_Wire_0[57], N263);
  xor keyGate_0_57(N300, keyinput57, keyinput_Wire_0[57]);
not NOT1_88 (N301, N288);
not NOT1_89 (N302, N289);
not NOT1_90 (N303, N290);
not NOT1_91 (N304, N291);
not NOT1_92 (N305, N292);
not NOT1_93 (N306, N293);
  not NOT1_94 (keyinput_Wire_0[58], N294);
  xnor keyGate_0_58(KeyNOTWire_0[24], keyinput58, keyinput_Wire_0[58]);
  not KeyNOTGate_0_24(N307, KeyNOTWire_0[24]);
not NOT1_95 (N308, N295);
not NOT1_96 (N309, N296);
not NOT1_97 (N319, N296);
not NOT1_98 (N329, N296);
xor XOR2_99 (N330, N309, N260);
  xor XOR2_100 (keyinput_Wire_0[59], N309, N264);
  xnor keyGate_0_59(KeyNOTWire_0[25], keyinput59, keyinput_Wire_0[59]);
  not KeyNOTGate_0_25(N331, KeyNOTWire_0[25]);
xor XOR2_101 (N332, N309, N267);
xor XOR2_102 (N333, N309, N270);
nand NAND2_103 (N334, N8, N319);
  xor XOR2_104 (keyinput_Wire_0[60], N309, N273);
  xor keyGate_0_60(N335, keyinput60, keyinput_Wire_0[60]);
nand NAND2_105 (N336, N319, N21);
xor XOR2_106 (N337, N309, N276);
nand NAND2_107 (N338, N319, N34);
xor XOR2_108 (N339, N309, N279);
nand NAND2_109 (N340, N319, N47);
xor XOR2_110 (N341, N309, N282);
nand NAND2_111 (N342, N319, N60);
xor XOR2_112 (N343, N309, N285);
nand NAND2_113 (N344, N319, N73);
nand NAND2_114 (N345, N319, N86);
nand NAND2_115 (N346, N319, N99);
nand NAND2_116 (N347, N319, N112);
nand NAND2_117 (N348, N330, N300);
  nand NAND2_118 (keyinput_Wire_0[61], N331, N301);
  xor keyGate_0_61(N349, keyinput61, keyinput_Wire_0[61]);
nand NAND2_119 (N350, N332, N302);
nand NAND2_120 (N351, N333, N303);
nand NAND2_121 (N352, N335, N304);
nand NAND2_122 (N353, N337, N305);
nand NAND2_123 (N354, N339, N306);
nand NAND2_124 (N355, N341, N307);
  nand NAND2_125 (keyinput_Wire_0[62], N343, N308);
  xor keyGate_0_62(N356, keyinput62, keyinput_Wire_0[62]);
and AND9_126 (N357, N348, N349, N350, N351, N352, N353, N354, N355, N356);
not NOT1_127 (N360, N357);
not NOT1_128 (N370, N357);
nand NAND2_129 (N371, N14, N360);
  nand NAND2_130 (keyinput_Wire_0[63], N360, N27);
  xnor keyGate_0_63(KeyNOTWire_0[26], keyinput63, keyinput_Wire_0[63]);
  not KeyNOTGate_0_26(N372, KeyNOTWire_0[26]);
nand NAND2_131 (N373, N360, N40);
nand NAND2_132 (N374, N360, N53);
nand NAND2_133 (N375, N360, N66);
nand NAND2_134 (N376, N360, N79);
nand NAND2_135 (N377, N360, N92);
nand NAND2_136 (N378, N360, N105);
nand NAND2_137 (N379, N360, N115);
nand NAND4_138 (N380, N4, N242, N334, N371);
nand NAND4_139 (N381, N246, N336, N372, N17);
nand NAND4_140 (N386, N250, N338, N373, N30);
nand NAND4_141 (N393, N254, N340, N374, N43);
nand NAND4_142 (N399, N255, N342, N375, N56);
nand NAND4_143 (N404, N256, N344, N376, N69);
nand NAND4_144 (N407, N257, N345, N377, N82);
nand NAND4_145 (N411, N258, N346, N378, N95);
nand NAND4_146 (N414, N259, N347, N379, N108);
not NOT1_147 (N415, N380);
and AND8_148 (N416, N381, N386, N393, N399, N404, N407, N411, N414);
not NOT1_149 (N417, N393);
not NOT1_150 (N418, N404);
not NOT1_151 (N419, N407);
not NOT1_152 (N420, N411);
nor NOR2_153 (N421, N415, N416);
nand NAND2_154 (N422, N386, N417);
nand NAND4_155 (N425, N386, N393, N418, N399);
nand NAND3_156 (N428, N399, N393, N419);
nand NAND4_157 (N429, N386, N393, N407, N420);
nand NAND4_158 (N430, N381, N386, N422, N399);
nand NAND4_159 (KeyWire_0_1, N381, N386, N425, N428);
  xor flip_it (N431, KeyWire_0_1, KeyWire_0_2 );
nand NAND4_160 (N432, N381, N422, N425, N429);

AntiSAT some_name( KeyWire_0_2, N108, N30, N43, N69, N60, N53, N11, N17, N89, N8, N99, N4, N24, N115, N27, N92, N66, N21, N73, N95, N76, N82, N50, N86, N37, N1, N47, N105, N40, N112, N102, N14, N56, N63, N34, N79, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135,
       keyinput136, keyinput137, keyinput138, keyinput139, keyinput140,
       keyinput141, keyinput142, keyinput143, keyinput144, keyinput145,
       keyinput146, keyinput147, keyinput148, keyinput149, keyinput150,
       keyinput151, keyinput152, keyinput153, keyinput154, keyinput155,
       keyinput156, keyinput157, keyinput158, keyinput159, keyinput160,
       keyinput161, keyinput162, keyinput163, keyinput164, keyinput165,
       keyinput166, keyinput167, keyinput168, keyinput169, keyinput170,
       keyinput171);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N108, N30, N43, N69, N60, N53, N11, N17, N89, N8, N99, N4, N24, N115, N27, N92, N66, N21, N73, N95, N76, N82, N50, N86, N37, N1, N47, N105, N40, N112, N102, N14, N56, N63, N34, N79, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135 ,
        keyinput136, keyinput137, keyinput138, keyinput139, keyinput140,
        keyinput141, keyinput142, keyinput143, keyinput144, keyinput145,
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150,
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155,
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160,
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165,
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170,
        keyinput171);

  input keyinput136, keyinput137, keyinput138, keyinput139, keyinput140;
  input keyinput141, keyinput142, keyinput143, keyinput144, keyinput145;
  input keyinput146, keyinput147, keyinput148, keyinput149, keyinput150;
  input keyinput151, keyinput152, keyinput153, keyinput154, keyinput155;
  input keyinput156, keyinput157, keyinput158, keyinput159, keyinput160;
  input keyinput161, keyinput162, keyinput163, keyinput164, keyinput165;
  input keyinput166, keyinput167, keyinput168, keyinput169, keyinput170;
  input keyinput171;

  wire [0:35] keyNTin_Wire_1;
  wire [0:15] KeyNOTWire_1;

  input N108, N30, N43, N69, N60, N53, N11, N17, N89, N8, N99, N4, N24, N115, N27, N92, N66, N21, N73, N95, N76, N82, N50, N86, N37, N1, N47, N105, N40, N112, N102, N14, N56, N63, N34, N79;
  input keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73 ;

  xnor KeyGate0 (newWire_0, N108, keyinput64);
  xor  KeyGate1 (newWire_1, N30, keyinput65);
  xnor KeyGate2 (keyNTin_Wire_1[0], N43, keyinput66);
  xor keyNTinGate_1_0(KeyNOTWire_1[0], keyinput136, keyNTin_Wire_1[0]);
  not KeyNOTGate_1_0(newWire_2, KeyNOTWire_1[0]);
  xor  KeyGate3 (newWire_3, N69, keyinput67);
  xnor KeyGate4 (keyNTin_Wire_1[1], N60, keyinput68);
  xor keyNTinGate_1_1(KeyNOTWire_1[1], keyinput137, keyNTin_Wire_1[1]);
  not KeyNOTGate_1_1(newWire_4, KeyNOTWire_1[1]);
  xnor KeyGate5 (keyNTin_Wire_1[2], N53, keyinput69);
  xnor keyNTinGate_1_2(newWire_5, keyinput138, keyNTin_Wire_1[2]);
  xor  KeyGate6 (keyNTin_Wire_1[3], N11, keyinput70);
  xnor keyNTinGate_1_3(KeyNOTWire_1[2], keyinput139, keyNTin_Wire_1[3]);
  not KeyNOTGate_1_2(newWire_6, KeyNOTWire_1[2]);
  xnor KeyGate7 (newWire_7, N17, keyinput71);
  xnor KeyGate8 (newWire_8, N89, keyinput72);
  xor  KeyGate9 (newWire_9, N8, keyinput73);
  xnor KeyGate10 (keyNTin_Wire_1[4], N99, keyinput74);
  xor keyNTinGate_1_4(newWire_10, keyinput140, keyNTin_Wire_1[4]);
  xor  KeyGate11 (newWire_11, N4, keyinput75);
  xor  KeyGate12 (keyNTin_Wire_1[5], N24, keyinput76);
  xor keyNTinGate_1_5(newWire_12, keyinput141, keyNTin_Wire_1[5]);
  xor  KeyGate13 (keyNTin_Wire_1[6], N115, keyinput77);
  xnor keyNTinGate_1_6(KeyNOTWire_1[3], keyinput142, keyNTin_Wire_1[6]);
  not KeyNOTGate_1_3(newWire_13, KeyNOTWire_1[3]);
  xor  KeyGate14 (newWire_14, N27, keyinput78);
  xor  KeyGate15 (newWire_15, N92, keyinput79);
  xnor KeyGate16 (newWire_16, N66, keyinput80);
  xnor KeyGate17 (keyNTin_Wire_1[7], N21, keyinput81);
  xnor keyNTinGate_1_7(KeyNOTWire_1[4], keyinput143, keyNTin_Wire_1[7]);
  not KeyNOTGate_1_4(newWire_17, KeyNOTWire_1[4]);
  xnor KeyGate18 (keyNTin_Wire_1[8], N73, keyinput82);
  xor keyNTinGate_1_8(newWire_18, keyinput144, keyNTin_Wire_1[8]);
  xnor KeyGate19 (newWire_19, N95, keyinput83);
  xor  KeyGate20 (newWire_20, N76, keyinput84);
  xor  KeyGate21 (keyNTin_Wire_1[9], N82, keyinput85);
  xnor keyNTinGate_1_9(newWire_21, keyinput145, keyNTin_Wire_1[9]);
  xnor KeyGate22 (keyNTin_Wire_1[10], N50, keyinput86);
  xnor keyNTinGate_1_10(newWire_22, keyinput146, keyNTin_Wire_1[10]);
  xnor KeyGate23 (newWire_23, N86, keyinput87);
  xnor KeyGate24 (newWire_24, N37, keyinput88);
  xor  KeyGate25 (newWire_25, N1, keyinput89);
  xor  KeyGate26 (newWire_26, N47, keyinput90);
  xnor KeyGate27 (newWire_27, N105, keyinput91);
  xor  KeyGate28 (newWire_28, N40, keyinput92);
  xor  KeyGate29 (newWire_29, N112, keyinput93);
  xor  KeyGate30 (keyNTin_Wire_1[11], N102, keyinput94);
  xnor keyNTinGate_1_11(newWire_30, keyinput147, keyNTin_Wire_1[11]);
  xor  KeyGate31 (newWire_31, N14, keyinput95);
  xnor KeyGate32 (keyNTin_Wire_1[12], N56, keyinput96);
  xnor keyNTinGate_1_12(newWire_32, keyinput148, keyNTin_Wire_1[12]);
  xnor KeyGate33 (newWire_33, N63, keyinput97);
  xnor KeyGate34 (newWire_34, N34, keyinput98);
  xor  KeyGate35 (newWire_35, N79, keyinput99);
  xnor KeyGate36 (newWire_36, N108, keyinput100);
  xnor KeyGate37 (keyNTin_Wire_1[13], N30, keyinput101);
  xor keyNTinGate_1_13(KeyNOTWire_1[5], keyinput149, keyNTin_Wire_1[13]);
  not KeyNOTGate_1_5(newWire_37, KeyNOTWire_1[5]);
  xor  KeyGate38 (keyNTin_Wire_1[14], N43, keyinput102);
  xnor keyNTinGate_1_14(newWire_38, keyinput150, keyNTin_Wire_1[14]);
  xor  KeyGate39 (keyNTin_Wire_1[15], N69, keyinput103);
  xor keyNTinGate_1_15(KeyNOTWire_1[6], keyinput151, keyNTin_Wire_1[15]);
  not KeyNOTGate_1_6(newWire_39, KeyNOTWire_1[6]);
  xnor KeyGate40 (keyNTin_Wire_1[16], N60, keyinput104);
  xnor keyNTinGate_1_16(KeyNOTWire_1[7], keyinput152, keyNTin_Wire_1[16]);
  not KeyNOTGate_1_7(newWire_40, KeyNOTWire_1[7]);
  xnor KeyGate41 (newWire_41, N53, keyinput105);
  xnor KeyGate42 (newWire_42, N11, keyinput106);
  xor  KeyGate43 (newWire_43, N17, keyinput107);
  xnor KeyGate44 (newWire_44, N89, keyinput108);
  xor  KeyGate45 (keyNTin_Wire_1[17], N8, keyinput109);
  xnor keyNTinGate_1_17(KeyNOTWire_1[8], keyinput153, keyNTin_Wire_1[17]);
  not KeyNOTGate_1_8(newWire_45, KeyNOTWire_1[8]);
  xor  KeyGate46 (keyNTin_Wire_1[18], N99, keyinput110);
  xnor keyNTinGate_1_18(newWire_46, keyinput154, keyNTin_Wire_1[18]);
  xnor KeyGate47 (keyNTin_Wire_1[19], N4, keyinput111);
  xor keyNTinGate_1_19(KeyNOTWire_1[9], keyinput155, keyNTin_Wire_1[19]);
  not KeyNOTGate_1_9(newWire_47, KeyNOTWire_1[9]);
  xor  KeyGate48 (newWire_48, N24, keyinput112);
  xnor KeyGate49 (newWire_49, N115, keyinput113);
  xor  KeyGate50 (newWire_50, N27, keyinput114);
  xor  KeyGate51 (newWire_51, N92, keyinput115);
  xnor KeyGate52 (newWire_52, N66, keyinput116);
  xor  KeyGate53 (keyNTin_Wire_1[20], N21, keyinput117);
  xor keyNTinGate_1_20(newWire_53, keyinput156, keyNTin_Wire_1[20]);
  xor  KeyGate54 (newWire_54, N73, keyinput118);
  xnor KeyGate55 (keyNTin_Wire_1[21], N95, keyinput119);
  xnor keyNTinGate_1_21(newWire_55, keyinput157, keyNTin_Wire_1[21]);
  xor  KeyGate56 (keyNTin_Wire_1[22], N76, keyinput120);
  xnor keyNTinGate_1_22(newWire_56, keyinput158, keyNTin_Wire_1[22]);
  xnor KeyGate57 (newWire_57, N82, keyinput121);
  xor  KeyGate58 (keyNTin_Wire_1[23], N50, keyinput122);
  xor keyNTinGate_1_23(newWire_58, keyinput159, keyNTin_Wire_1[23]);
  xnor KeyGate59 (keyNTin_Wire_1[24], N86, keyinput123);
  xor keyNTinGate_1_24(newWire_59, keyinput160, keyNTin_Wire_1[24]);
  xnor KeyGate60 (keyNTin_Wire_1[25], N37, keyinput124);
  xnor keyNTinGate_1_25(newWire_60, keyinput161, keyNTin_Wire_1[25]);
  xnor KeyGate61 (keyNTin_Wire_1[26], N1, keyinput125);
  xor keyNTinGate_1_26(newWire_61, keyinput162, keyNTin_Wire_1[26]);
  xnor KeyGate62 (newWire_62, N47, keyinput126);
  xor  KeyGate63 (keyNTin_Wire_1[27], N105, keyinput127);
  xnor keyNTinGate_1_27(newWire_63, keyinput163, keyNTin_Wire_1[27]);
  xor  KeyGate64 (keyNTin_Wire_1[28], N40, keyinput128);
  xor keyNTinGate_1_28(newWire_64, keyinput164, keyNTin_Wire_1[28]);
  xor  KeyGate65 (keyNTin_Wire_1[29], N112, keyinput129);
  xor keyNTinGate_1_29(KeyNOTWire_1[10], keyinput165, keyNTin_Wire_1[29]);
  not KeyNOTGate_1_10(newWire_65, KeyNOTWire_1[10]);
  xnor KeyGate66 (newWire_66, N102, keyinput130);
  xnor KeyGate67 (keyNTin_Wire_1[30], N14, keyinput131);
  xor keyNTinGate_1_30(KeyNOTWire_1[11], keyinput166, keyNTin_Wire_1[30]);
  not KeyNOTGate_1_11(newWire_67, KeyNOTWire_1[11]);
  xnor KeyGate68 (keyNTin_Wire_1[31], N56, keyinput132);
  xor keyNTinGate_1_31(newWire_68, keyinput167, keyNTin_Wire_1[31]);
  xor  KeyGate69 (newWire_69, N63, keyinput133);
  xor  KeyGate70 (keyNTin_Wire_1[32], N34, keyinput134);
  xor keyNTinGate_1_32(KeyNOTWire_1[12], keyinput168, keyNTin_Wire_1[32]);
  not KeyNOTGate_1_12(newWire_70, KeyNOTWire_1[12]);
  xor  KeyGate71 (keyNTin_Wire_1[33], N79, keyinput135);
  xor keyNTinGate_1_33(KeyNOTWire_1[13], keyinput169, keyNTin_Wire_1[33]);
  not KeyNOTGate_1_13(newWire_71, KeyNOTWire_1[13]);
  and some_function (keyNTin_Wire_1[34], newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35 );
  xor keyNTinGate_1_34(KeyNOTWire_1[14], keyinput170, keyNTin_Wire_1[34]);
  not KeyNOTGate_1_14(newWire_72, KeyNOTWire_1[14]);
  nand compl_function (keyNTin_Wire_1[35], newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71);
  xor keyNTinGate_1_35(KeyNOTWire_1[15], keyinput171, keyNTin_Wire_1[35]);
  not KeyNOTGate_1_15(newWire_73, KeyNOTWire_1[15]);
  and finalAND (KeyWire_0_2, newWire_72, newWire_73);

endmodule /* AntiSAT */
