`timescale 1ns / 1ps
// Verilog
// c1908
// Ninputs 33
// Noutputs 25
// NtotalGates 880
// NOT1 277
// NAND2 347
// BUFF1 162
// AND2 30
// AND3 12
// NAND4 2
// NAND3 1
// NAND8 3
// AND4 2
// NAND5 24
// AND5 16
// AND8 3
// NOR2 1

module top (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
                  N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899,
        keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4,
        keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9,
        keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14,
        keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19,
        keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24,
        keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29,
        keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34,
        keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39,
        keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44,
        keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49,
        keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54,
        keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59,
        keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64,
        keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69,
        keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74,
        keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79,
        keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84,
        keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89,
        keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94,
        keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99,
        keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104,
        keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109,
        keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114,
        keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119,
        keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124,
        keyIn_0_125, keyIn_0_126, keyIn_0_127);

  input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4;
  input keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9;
  input keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14;
  input keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19;
  input keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24;
  input keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29;
  input keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34;
  input keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39;
  input keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44;
  input keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49;
  input keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54;
  input keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59;
  input keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64;
  input keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69;
  input keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74;
  input keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79;
  input keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84;
  input keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89;
  input keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94;
  input keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99;
  input keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104;
  input keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109;
  input keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114;
  input keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119;
  input keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124;
  input keyIn_0_125, keyIn_0_126, keyIn_0_127;

  wire [0:127] KeyWire_0;
  wire [0:71] KeyNOTWire_0;

input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;

output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;

wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898;

not NOT1_1 (N190, N1);
not NOT1_2 (N194, N4);
not NOT1_3 (N197, N7);
not NOT1_4 (N201, N10);
not NOT1_5 (N206, N13);
not NOT1_6 (N209, N16);
not NOT1_7 (N212, N19);
not NOT1_8 (N216, N22);
not NOT1_9 (N220, N25);
not NOT1_10 (N225, N28);
not NOT1_11 (N229, N31);
not NOT1_12 (N232, N34);
not NOT1_13 (N235, N37);
not NOT1_14 (N239, N40);
not NOT1_15 (N243, N43);
not NOT1_16 (N247, N46);
nand NAND2_17 (N251, N63, N88);
nand NAND2_18 (N252, N66, N91);
not NOT1_19 (N253, N72);
not NOT1_20 (N256, N72);
buf BUFF1_21 (N257, N69);
buf BUFF1_22 (N260, N69);
not NOT1_23 (N263, N76);
not NOT1_24 (N266, N79);
not NOT1_25 (N269, N82);
not NOT1_26 (N272, N85);
not NOT1_27 (N275, N104);
not NOT1_28 (N276, N104);
  not NOT1_29 (KeyWire_0[0], N88);
  xor KeyGate_0_0(N277, keyIn_0_0, KeyWire_0[0]);
  not NOT1_30 (KeyWire_0[1], N91);
  xnor KeyGate_0_1(KeyNOTWire_0[0], keyIn_0_1, KeyWire_0[1]);
  not KeyNOTGate_0_0(N280, KeyNOTWire_0[0]);
buf BUFF1_31 (N283, N94);
not NOT1_32 (N290, N94);
buf BUFF1_33 (N297, N94);
not NOT1_34 (N300, N94);
buf BUFF1_35 (N303, N99);
not NOT1_36 (N306, N99);
not NOT1_37 (N313, N99);
buf BUFF1_38 (N316, N104);
not NOT1_39 (N319, N104);
buf BUFF1_40 (N326, N104);
buf BUFF1_41 (N331, N104);
  not NOT1_42 (KeyWire_0[2], N104);
  xnor KeyGate_0_2(KeyNOTWire_0[1], keyIn_0_2, KeyWire_0[2]);
  not KeyNOTGate_0_1(N338, KeyNOTWire_0[1]);
buf BUFF1_43 (N343, N1);
buf BUFF1_44 (N346, N4);
buf BUFF1_45 (N349, N7);
buf BUFF1_46 (N352, N10);
buf BUFF1_47 (N355, N13);
buf BUFF1_48 (N358, N16);
buf BUFF1_49 (N361, N19);
buf BUFF1_50 (N364, N22);
buf BUFF1_51 (N367, N25);
buf BUFF1_52 (N370, N28);
buf BUFF1_53 (N373, N31);
buf BUFF1_54 (N376, N34);
buf BUFF1_55 (N379, N37);
buf BUFF1_56 (N382, N40);
buf BUFF1_57 (N385, N43);
buf BUFF1_58 (N388, N46);
not NOT1_59 (N534, N343);
not NOT1_60 (N535, N346);
not NOT1_61 (N536, N349);
not NOT1_62 (N537, N352);
not NOT1_63 (N538, N355);
not NOT1_64 (N539, N358);
not NOT1_65 (N540, N361);
not NOT1_66 (N541, N364);
not NOT1_67 (N542, N367);
not NOT1_68 (N543, N370);
not NOT1_69 (N544, N373);
not NOT1_70 (N545, N376);
not NOT1_71 (N546, N379);
not NOT1_72 (N547, N382);
not NOT1_73 (N548, N385);
not NOT1_74 (N549, N388);
nand NAND2_75 (N550, N306, N331);
nand NAND2_76 (N551, N306, N331);
nand NAND2_77 (N552, N306, N331);
nand NAND2_78 (N553, N306, N331);
nand NAND2_79 (N554, N306, N331);
nand NAND2_80 (N555, N306, N331);
buf BUFF1_81 (N556, N190);
buf BUFF1_82 (N559, N194);
buf BUFF1_83 (N562, N206);
buf BUFF1_84 (N565, N209);
buf BUFF1_85 (N568, N225);
buf BUFF1_86 (N571, N243);
and AND2_87 (N574, N63, N319);
buf BUFF1_88 (N577, N220);
buf BUFF1_89 (N580, N229);
buf BUFF1_90 (N583, N232);
and AND2_91 (N586, N66, N319);
buf BUFF1_92 (N589, N239);
and AND3_93 (N592, N49, N253, N319);
buf BUFF1_94 (N595, N247);
buf BUFF1_95 (N598, N239);
nand NAND2_96 (N601, N326, N277);
nand NAND2_97 (N602, N326, N280);
  nand NAND2_98 (KeyWire_0[3], N260, N72);
  xnor KeyGate_0_3(KeyNOTWire_0[2], keyIn_0_3, KeyWire_0[3]);
  not KeyNOTGate_0_2(N603, KeyNOTWire_0[2]);
nand NAND2_99 (N608, N260, N300);
nand NAND2_100 (N612, N256, N300);
buf BUFF1_101 (N616, N201);
buf BUFF1_102 (N619, N216);
buf BUFF1_103 (N622, N220);
buf BUFF1_104 (N625, N239);
buf BUFF1_105 (N628, N190);
buf BUFF1_106 (N631, N190);
buf BUFF1_107 (N634, N194);
buf BUFF1_108 (N637, N229);
buf BUFF1_109 (N640, N197);
and AND3_110 (N643, N56, N257, N319);
buf BUFF1_111 (N646, N232);
buf BUFF1_112 (N649, N201);
buf BUFF1_113 (N652, N235);
and AND3_114 (N655, N60, N257, N319);
buf BUFF1_115 (N658, N263);
buf BUFF1_116 (N661, N263);
buf BUFF1_117 (N664, N266);
buf BUFF1_118 (N667, N266);
buf BUFF1_119 (N670, N269);
buf BUFF1_120 (N673, N269);
buf BUFF1_121 (N676, N272);
buf BUFF1_122 (N679, N272);
and AND2_123 (N682, N251, N316);
and AND2_124 (N685, N252, N316);
buf BUFF1_125 (N688, N197);
buf BUFF1_126 (N691, N197);
buf BUFF1_127 (N694, N212);
buf BUFF1_128 (N697, N212);
buf BUFF1_129 (N700, N247);
buf BUFF1_130 (N703, N247);
buf BUFF1_131 (N706, N235);
buf BUFF1_132 (N709, N235);
buf BUFF1_133 (N712, N201);
buf BUFF1_134 (N715, N201);
buf BUFF1_135 (N718, N206);
buf BUFF1_136 (N721, N216);
and AND3_137 (N724, N53, N253, N319);
buf BUFF1_138 (N727, N243);
buf BUFF1_139 (N730, N220);
buf BUFF1_140 (N733, N220);
buf BUFF1_141 (N736, N209);
buf BUFF1_142 (N739, N216);
buf BUFF1_143 (N742, N225);
buf BUFF1_144 (N745, N243);
buf BUFF1_145 (N748, N212);
buf BUFF1_146 (N751, N225);
not NOT1_147 (N886, N682);
not NOT1_148 (N887, N685);
not NOT1_149 (N888, N616);
not NOT1_150 (N889, N619);
not NOT1_151 (N890, N622);
  not NOT1_152 (KeyWire_0[4], N625);
  xnor KeyGate_0_4(KeyNOTWire_0[3], keyIn_0_4, KeyWire_0[4]);
  not KeyNOTGate_0_3(N891, KeyNOTWire_0[3]);
not NOT1_153 (N892, N631);
not NOT1_154 (N893, N643);
not NOT1_155 (N894, N649);
not NOT1_156 (N895, N652);
not NOT1_157 (N896, N655);
  and AND2_158 (KeyWire_0[5], N49, N612);
  xor KeyGate_0_5(N897, keyIn_0_5, KeyWire_0[5]);
and AND2_159 (N898, N56, N608);
nand NAND2_160 (N899, N53, N612);
nand NAND2_161 (N903, N60, N608);
nand NAND2_162 (N907, N49, N612);
nand NAND2_163 (N910, N56, N608);
not NOT1_164 (N913, N661);
  not NOT1_165 (KeyWire_0[6], N658);
  xor KeyGate_0_6(KeyNOTWire_0[4], keyIn_0_6, KeyWire_0[6]);
  not KeyNOTGate_0_4(N914, KeyNOTWire_0[4]);
not NOT1_166 (N915, N667);
  not NOT1_167 (KeyWire_0[7], N664);
  xnor KeyGate_0_7(N916, keyIn_0_7, KeyWire_0[7]);
not NOT1_168 (N917, N673);
  not NOT1_169 (KeyWire_0[8], N670);
  xnor KeyGate_0_8(N918, keyIn_0_8, KeyWire_0[8]);
not NOT1_170 (N919, N679);
  not NOT1_171 (KeyWire_0[9], N676);
  xor KeyGate_0_9(KeyNOTWire_0[5], keyIn_0_9, KeyWire_0[9]);
  not KeyNOTGate_0_5(N920, KeyNOTWire_0[5]);
  nand NAND4_172 (KeyWire_0[10], N277, N297, N326, N603);
  xnor KeyGate_0_10(KeyNOTWire_0[6], keyIn_0_10, KeyWire_0[10]);
  not KeyNOTGate_0_6(N921, KeyNOTWire_0[6]);
  nand NAND4_173 (KeyWire_0[11], N280, N297, N326, N603);
  xor KeyGate_0_11(KeyNOTWire_0[7], keyIn_0_11, KeyWire_0[11]);
  not KeyNOTGate_0_7(N922, KeyNOTWire_0[7]);
  nand NAND3_174 (KeyWire_0[12], N303, N338, N603);
  xnor KeyGate_0_12(N923, keyIn_0_12, KeyWire_0[12]);
and AND3_175 (N926, N303, N338, N603);
buf BUFF1_176 (N935, N556);
not NOT1_177 (N938, N688);
buf BUFF1_178 (N939, N556);
not NOT1_179 (N942, N691);
buf BUFF1_180 (N943, N562);
not NOT1_181 (N946, N694);
buf BUFF1_182 (N947, N562);
  not NOT1_183 (KeyWire_0[13], N697);
  xnor KeyGate_0_13(N950, keyIn_0_13, KeyWire_0[13]);
buf BUFF1_184 (N951, N568);
not NOT1_185 (N954, N700);
buf BUFF1_186 (N955, N568);
not NOT1_187 (N958, N703);
buf BUFF1_188 (N959, N574);
buf BUFF1_189 (N962, N574);
buf BUFF1_190 (N965, N580);
not NOT1_191 (N968, N706);
buf BUFF1_192 (N969, N580);
not NOT1_193 (N972, N709);
buf BUFF1_194 (N973, N586);
not NOT1_195 (N976, N712);
buf BUFF1_196 (N977, N586);
not NOT1_197 (N980, N715);
buf BUFF1_198 (N981, N592);
not NOT1_199 (N984, N628);
buf BUFF1_200 (N985, N592);
not NOT1_201 (N988, N718);
not NOT1_202 (N989, N721);
not NOT1_203 (N990, N634);
not NOT1_204 (N991, N724);
not NOT1_205 (N992, N727);
not NOT1_206 (N993, N637);
buf BUFF1_207 (N994, N595);
not NOT1_208 (N997, N730);
buf BUFF1_209 (N998, N595);
not NOT1_210 (N1001, N733);
not NOT1_211 (N1002, N736);
not NOT1_212 (N1003, N739);
not NOT1_213 (N1004, N640);
not NOT1_214 (N1005, N742);
not NOT1_215 (N1006, N745);
not NOT1_216 (N1007, N646);
not NOT1_217 (N1008, N748);
not NOT1_218 (N1009, N751);
buf BUFF1_219 (N1010, N559);
buf BUFF1_220 (N1013, N559);
buf BUFF1_221 (N1016, N565);
buf BUFF1_222 (N1019, N565);
buf BUFF1_223 (N1022, N571);
buf BUFF1_224 (N1025, N571);
buf BUFF1_225 (N1028, N577);
buf BUFF1_226 (N1031, N577);
buf BUFF1_227 (N1034, N583);
buf BUFF1_228 (N1037, N583);
buf BUFF1_229 (N1040, N589);
buf BUFF1_230 (N1043, N589);
buf BUFF1_231 (N1046, N598);
buf BUFF1_232 (N1049, N598);
nand NAND2_233 (N1054, N619, N888);
nand NAND2_234 (N1055, N616, N889);
nand NAND2_235 (N1063, N625, N890);
nand NAND2_236 (N1064, N622, N891);
nand NAND2_237 (N1067, N655, N895);
nand NAND2_238 (N1068, N652, N896);
nand NAND2_239 (N1119, N721, N988);
nand NAND2_240 (N1120, N718, N989);
nand NAND2_241 (N1121, N727, N991);
nand NAND2_242 (N1122, N724, N992);
nand NAND2_243 (N1128, N739, N1002);
nand NAND2_244 (N1129, N736, N1003);
nand NAND2_245 (N1130, N745, N1005);
nand NAND2_246 (N1131, N742, N1006);
nand NAND2_247 (N1132, N751, N1008);
nand NAND2_248 (N1133, N748, N1009);
not NOT1_249 (N1148, N939);
  not NOT1_250 (KeyWire_0[14], N935);
  xnor KeyGate_0_14(N1149, keyIn_0_14, KeyWire_0[14]);
nand NAND2_251 (N1150, N1054, N1055);
not NOT1_252 (N1151, N943);
not NOT1_253 (N1152, N947);
not NOT1_254 (N1153, N955);
not NOT1_255 (N1154, N951);
not NOT1_256 (N1155, N962);
not NOT1_257 (N1156, N969);
not NOT1_258 (N1157, N977);
nand NAND2_259 (N1158, N1063, N1064);
not NOT1_260 (N1159, N985);
nand NAND2_261 (N1160, N985, N892);
not NOT1_262 (N1161, N998);
nand NAND2_263 (N1162, N1067, N1068);
not NOT1_264 (N1163, N899);
buf BUFF1_265 (N1164, N899);
not NOT1_266 (N1167, N903);
buf BUFF1_267 (N1168, N903);
  nand NAND2_268 (KeyWire_0[15], N921, N923);
  xnor KeyGate_0_15(KeyNOTWire_0[8], keyIn_0_15, KeyWire_0[15]);
  not KeyNOTGate_0_8(N1171, KeyNOTWire_0[8]);
  nand NAND2_269 (KeyWire_0[16], N922, N923);
  xor KeyGate_0_16(N1188, keyIn_0_16, KeyWire_0[16]);
not NOT1_270 (N1205, N1010);
nand NAND2_271 (N1206, N1010, N938);
not NOT1_272 (N1207, N1013);
nand NAND2_273 (N1208, N1013, N942);
not NOT1_274 (N1209, N1016);
nand NAND2_275 (N1210, N1016, N946);
not NOT1_276 (N1211, N1019);
nand NAND2_277 (N1212, N1019, N950);
not NOT1_278 (N1213, N1022);
nand NAND2_279 (N1214, N1022, N954);
not NOT1_280 (N1215, N1025);
nand NAND2_281 (N1216, N1025, N958);
not NOT1_282 (N1217, N1028);
not NOT1_283 (N1218, N959);
not NOT1_284 (N1219, N1031);
not NOT1_285 (N1220, N1034);
nand NAND2_286 (N1221, N1034, N968);
not NOT1_287 (N1222, N965);
not NOT1_288 (N1223, N1037);
nand NAND2_289 (N1224, N1037, N972);
not NOT1_290 (N1225, N1040);
nand NAND2_291 (N1226, N1040, N976);
not NOT1_292 (N1227, N973);
not NOT1_293 (N1228, N1043);
nand NAND2_294 (N1229, N1043, N980);
not NOT1_295 (N1230, N981);
nand NAND2_296 (N1231, N981, N984);
nand NAND2_297 (N1232, N1119, N1120);
nand NAND2_298 (N1235, N1121, N1122);
not NOT1_299 (N1238, N1046);
nand NAND2_300 (N1239, N1046, N997);
not NOT1_301 (N1240, N994);
not NOT1_302 (N1241, N1049);
nand NAND2_303 (N1242, N1049, N1001);
nand NAND2_304 (N1243, N1128, N1129);
nand NAND2_305 (N1246, N1130, N1131);
nand NAND2_306 (N1249, N1132, N1133);
buf BUFF1_307 (N1252, N907);
buf BUFF1_308 (N1255, N907);
buf BUFF1_309 (N1258, N910);
buf BUFF1_310 (N1261, N910);
not NOT1_311 (N1264, N1150);
nand NAND2_312 (N1267, N631, N1159);
nand NAND2_313 (N1309, N688, N1205);
nand NAND2_314 (N1310, N691, N1207);
nand NAND2_315 (N1311, N694, N1209);
nand NAND2_316 (N1312, N697, N1211);
nand NAND2_317 (N1313, N700, N1213);
nand NAND2_318 (N1314, N703, N1215);
nand NAND2_319 (N1315, N706, N1220);
nand NAND2_320 (N1316, N709, N1223);
nand NAND2_321 (N1317, N712, N1225);
nand NAND2_322 (N1318, N715, N1228);
not NOT1_323 (N1319, N1158);
nand NAND2_324 (N1322, N628, N1230);
nand NAND2_325 (N1327, N730, N1238);
nand NAND2_326 (N1328, N733, N1241);
not NOT1_327 (N1334, N1162);
nand NAND2_328 (N1344, N1267, N1160);
nand NAND2_329 (N1345, N1249, N894);
not NOT1_330 (N1346, N1249);
not NOT1_331 (N1348, N1255);
  not NOT1_332 (KeyWire_0[17], N1252);
  xor KeyGate_0_17(KeyNOTWire_0[9], keyIn_0_17, KeyWire_0[17]);
  not KeyNOTGate_0_9(N1349, KeyNOTWire_0[9]);
not NOT1_333 (N1350, N1261);
  not NOT1_334 (KeyWire_0[18], N1258);
  xor KeyGate_0_18(N1351, keyIn_0_18, KeyWire_0[18]);
nand NAND2_335 (N1352, N1309, N1206);
nand NAND2_336 (N1355, N1310, N1208);
nand NAND2_337 (N1358, N1311, N1210);
  nand NAND2_338 (KeyWire_0[19], N1312, N1212);
  xor KeyGate_0_19(KeyNOTWire_0[10], keyIn_0_19, KeyWire_0[19]);
  not KeyNOTGate_0_10(N1361, KeyNOTWire_0[10]);
nand NAND2_339 (N1364, N1313, N1214);
nand NAND2_340 (N1367, N1314, N1216);
nand NAND2_341 (N1370, N1315, N1221);
nand NAND2_342 (N1373, N1316, N1224);
nand NAND2_343 (N1376, N1317, N1226);
nand NAND2_344 (N1379, N1318, N1229);
nand NAND2_345 (N1383, N1322, N1231);
not NOT1_346 (N1386, N1232);
nand NAND2_347 (N1387, N1232, N990);
not NOT1_348 (N1388, N1235);
nand NAND2_349 (N1389, N1235, N993);
nand NAND2_350 (N1390, N1327, N1239);
nand NAND2_351 (N1393, N1328, N1242);
not NOT1_352 (N1396, N1243);
nand NAND2_353 (N1397, N1243, N1004);
not NOT1_354 (N1398, N1246);
nand NAND2_355 (N1399, N1246, N1007);
not NOT1_356 (N1409, N1319);
nand NAND2_357 (N1412, N649, N1346);
not NOT1_358 (N1413, N1334);
buf BUFF1_359 (N1416, N1264);
buf BUFF1_360 (N1419, N1264);
nand NAND2_361 (N1433, N634, N1386);
nand NAND2_362 (N1434, N637, N1388);
nand NAND2_363 (N1438, N640, N1396);
nand NAND2_364 (N1439, N646, N1398);
not NOT1_365 (N1440, N1344);
nand NAND2_366 (N1443, N1355, N1148);
not NOT1_367 (N1444, N1355);
nand NAND2_368 (N1445, N1352, N1149);
not NOT1_369 (N1446, N1352);
nand NAND2_370 (N1447, N1358, N1151);
not NOT1_371 (N1448, N1358);
nand NAND2_372 (N1451, N1361, N1152);
not NOT1_373 (N1452, N1361);
nand NAND2_374 (N1453, N1367, N1153);
not NOT1_375 (N1454, N1367);
nand NAND2_376 (N1455, N1364, N1154);
not NOT1_377 (N1456, N1364);
nand NAND2_378 (N1457, N1373, N1156);
not NOT1_379 (N1458, N1373);
nand NAND2_380 (N1459, N1379, N1157);
not NOT1_381 (N1460, N1379);
not NOT1_382 (N1461, N1383);
nand NAND2_383 (N1462, N1393, N1161);
not NOT1_384 (N1463, N1393);
nand NAND2_385 (N1464, N1345, N1412);
not NOT1_386 (N1468, N1370);
nand NAND2_387 (N1469, N1370, N1222);
not NOT1_388 (N1470, N1376);
nand NAND2_389 (N1471, N1376, N1227);
nand NAND2_390 (N1472, N1387, N1433);
not NOT1_391 (N1475, N1390);
nand NAND2_392 (N1476, N1390, N1240);
nand NAND2_393 (N1478, N1389, N1434);
nand NAND2_394 (N1481, N1399, N1439);
nand NAND2_395 (N1484, N1397, N1438);
nand NAND2_396 (N1487, N939, N1444);
nand NAND2_397 (N1488, N935, N1446);
nand NAND2_398 (N1489, N943, N1448);
not NOT1_399 (N1490, N1419);
not NOT1_400 (N1491, N1416);
nand NAND2_401 (N1492, N947, N1452);
nand NAND2_402 (N1493, N955, N1454);
nand NAND2_403 (N1494, N951, N1456);
nand NAND2_404 (N1495, N969, N1458);
nand NAND2_405 (N1496, N977, N1460);
nand NAND2_406 (N1498, N998, N1463);
not NOT1_407 (N1499, N1440);
nand NAND2_408 (N1500, N965, N1468);
nand NAND2_409 (N1501, N973, N1470);
nand NAND2_410 (N1504, N994, N1475);
not NOT1_411 (N1510, N1464);
nand NAND2_412 (N1513, N1443, N1487);
nand NAND2_413 (N1514, N1445, N1488);
nand NAND2_414 (N1517, N1447, N1489);
nand NAND2_415 (N1520, N1451, N1492);
nand NAND2_416 (N1521, N1453, N1493);
nand NAND2_417 (N1522, N1455, N1494);
nand NAND2_418 (N1526, N1457, N1495);
nand NAND2_419 (N1527, N1459, N1496);
not NOT1_420 (N1528, N1472);
nand NAND2_421 (N1529, N1462, N1498);
  not NOT1_422 (KeyWire_0[20], N1478);
  xnor KeyGate_0_20(N1530, keyIn_0_20, KeyWire_0[20]);
not NOT1_423 (N1531, N1481);
not NOT1_424 (N1532, N1484);
nand NAND2_425 (N1534, N1471, N1501);
nand NAND2_426 (N1537, N1469, N1500);
nand NAND2_427 (N1540, N1476, N1504);
not NOT1_428 (N1546, N1513);
not NOT1_429 (N1554, N1521);
not NOT1_430 (N1557, N1526);
not NOT1_431 (N1561, N1520);
  nand NAND2_432 (KeyWire_0[21], N1484, N1531);
  xnor KeyGate_0_21(KeyNOTWire_0[11], keyIn_0_21, KeyWire_0[21]);
  not KeyNOTGate_0_11(N1567, KeyNOTWire_0[11]);
nand NAND2_433 (N1568, N1481, N1532);
  not NOT1_434 (KeyWire_0[22], N1510);
  xnor KeyGate_0_22(KeyNOTWire_0[12], keyIn_0_22, KeyWire_0[22]);
  not KeyNOTGate_0_12(N1569, KeyNOTWire_0[12]);
not NOT1_435 (N1571, N1527);
not NOT1_436 (N1576, N1529);
buf BUFF1_437 (N1588, N1522);
not NOT1_438 (N1591, N1534);
not NOT1_439 (N1593, N1537);
nand NAND2_440 (N1594, N1540, N1530);
not NOT1_441 (N1595, N1540);
nand NAND2_442 (N1596, N1567, N1568);
buf BUFF1_443 (N1600, N1517);
buf BUFF1_444 (N1603, N1517);
buf BUFF1_445 (N1606, N1522);
buf BUFF1_446 (N1609, N1522);
buf BUFF1_447 (N1612, N1514);
buf BUFF1_448 (N1615, N1514);
buf BUFF1_449 (N1620, N1557);
buf BUFF1_450 (N1623, N1554);
not NOT1_451 (N1635, N1571);
nand NAND2_452 (N1636, N1478, N1595);
nand NAND2_453 (N1638, N1576, N1569);
not NOT1_454 (N1639, N1576);
buf BUFF1_455 (N1640, N1561);
buf BUFF1_456 (N1643, N1561);
buf BUFF1_457 (N1647, N1546);
buf BUFF1_458 (N1651, N1546);
buf BUFF1_459 (N1658, N1554);
buf BUFF1_460 (N1661, N1557);
buf BUFF1_461 (N1664, N1557);
nand NAND2_462 (N1671, N1596, N893);
not NOT1_463 (N1672, N1596);
not NOT1_464 (N1675, N1600);
not NOT1_465 (N1677, N1603);
nand NAND2_466 (N1678, N1606, N1217);
not NOT1_467 (N1679, N1606);
nand NAND2_468 (N1680, N1609, N1219);
not NOT1_469 (N1681, N1609);
not NOT1_470 (N1682, N1612);
not NOT1_471 (N1683, N1615);
nand NAND2_472 (N1685, N1594, N1636);
nand NAND2_473 (N1688, N1510, N1639);
buf BUFF1_474 (N1697, N1588);
buf BUFF1_475 (N1701, N1588);
nand NAND2_476 (N1706, N643, N1672);
not NOT1_477 (N1707, N1643);
nand NAND2_478 (N1708, N1647, N1675);
not NOT1_479 (N1709, N1647);
nand NAND2_480 (N1710, N1651, N1677);
not NOT1_481 (N1711, N1651);
nand NAND2_482 (N1712, N1028, N1679);
nand NAND2_483 (N1713, N1031, N1681);
buf BUFF1_484 (N1714, N1620);
buf BUFF1_485 (N1717, N1620);
nand NAND2_486 (N1720, N1658, N1593);
not NOT1_487 (N1721, N1658);
nand NAND2_488 (N1723, N1638, N1688);
not NOT1_489 (N1727, N1661);
not NOT1_490 (N1728, N1640);
not NOT1_491 (N1730, N1664);
buf BUFF1_492 (N1731, N1623);
buf BUFF1_493 (N1734, N1623);
nand NAND2_494 (N1740, N1685, N1528);
not NOT1_495 (N1741, N1685);
nand NAND2_496 (N1742, N1671, N1706);
nand NAND2_497 (N1746, N1600, N1709);
nand NAND2_498 (N1747, N1603, N1711);
nand NAND2_499 (N1748, N1678, N1712);
nand NAND2_500 (N1751, N1680, N1713);
nand NAND2_501 (N1759, N1537, N1721);
not NOT1_502 (N1761, N1697);
nand NAND2_503 (N1762, N1697, N1727);
not NOT1_504 (N1763, N1701);
nand NAND2_505 (N1764, N1701, N1730);
not NOT1_506 (N1768, N1717);
nand NAND2_507 (N1769, N1472, N1741);
nand NAND2_508 (N1772, N1723, N1413);
not NOT1_509 (N1773, N1723);
nand NAND2_510 (N1774, N1708, N1746);
nand NAND2_511 (N1777, N1710, N1747);
not NOT1_512 (N1783, N1731);
nand NAND2_513 (N1784, N1731, N1682);
not NOT1_514 (N1785, N1714);
not NOT1_515 (N1786, N1734);
nand NAND2_516 (N1787, N1734, N1683);
nand NAND2_517 (N1788, N1720, N1759);
nand NAND2_518 (N1791, N1661, N1761);
nand NAND2_519 (N1792, N1664, N1763);
nand NAND2_520 (N1795, N1751, N1155);
not NOT1_521 (N1796, N1751);
nand NAND2_522 (N1798, N1740, N1769);
  nand NAND2_523 (KeyWire_0[23], N1334, N1773);
  xor KeyGate_0_23(KeyNOTWire_0[13], keyIn_0_23, KeyWire_0[23]);
  not KeyNOTGate_0_13(N1801, KeyNOTWire_0[13]);
nand NAND2_524 (N1802, N1742, N290);
not NOT1_525 (N1807, N1748);
nand NAND2_526 (N1808, N1748, N1218);
nand NAND2_527 (N1809, N1612, N1783);
nand NAND2_528 (N1810, N1615, N1786);
nand NAND2_529 (N1812, N1791, N1762);
nand NAND2_530 (N1815, N1792, N1764);
buf BUFF1_531 (N1818, N1742);
nand NAND2_532 (N1821, N1777, N1490);
not NOT1_533 (N1822, N1777);
nand NAND2_534 (N1823, N1774, N1491);
not NOT1_535 (N1824, N1774);
nand NAND2_536 (N1825, N962, N1796);
nand NAND2_537 (N1826, N1788, N1409);
not NOT1_538 (N1827, N1788);
nand NAND2_539 (N1830, N1772, N1801);
nand NAND2_540 (N1837, N959, N1807);
nand NAND2_541 (N1838, N1809, N1784);
nand NAND2_542 (N1841, N1810, N1787);
nand NAND2_543 (N1848, N1419, N1822);
nand NAND2_544 (N1849, N1416, N1824);
nand NAND2_545 (N1850, N1795, N1825);
nand NAND2_546 (N1852, N1319, N1827);
nand NAND2_547 (N1855, N1815, N1707);
not NOT1_548 (N1856, N1815);
not NOT1_549 (N1857, N1818);
nand NAND2_550 (N1858, N1798, N290);
not NOT1_551 (N1864, N1812);
nand NAND2_552 (N1865, N1812, N1728);
buf BUFF1_553 (N1866, N1798);
buf BUFF1_554 (N1869, N1802);
buf BUFF1_555 (N1872, N1802);
nand NAND2_556 (N1875, N1808, N1837);
nand NAND2_557 (N1878, N1821, N1848);
nand NAND2_558 (N1879, N1823, N1849);
nand NAND2_559 (N1882, N1841, N1768);
not NOT1_560 (N1883, N1841);
nand NAND2_561 (N1884, N1826, N1852);
nand NAND2_562 (N1885, N1643, N1856);
nand NAND2_563 (N1889, N1830, N290);
not NOT1_564 (N1895, N1838);
nand NAND2_565 (N1896, N1838, N1785);
nand NAND2_566 (N1897, N1640, N1864);
not NOT1_567 (N1898, N1850);
buf BUFF1_568 (N1902, N1830);
not NOT1_569 (N1910, N1878);
nand NAND2_570 (N1911, N1717, N1883);
not NOT1_571 (N1912, N1884);
nand NAND2_572 (N1913, N1855, N1885);
not NOT1_573 (N1915, N1866);
nand NAND2_574 (N1919, N1872, N919);
not NOT1_575 (N1920, N1872);
  nand NAND2_576 (KeyWire_0[24], N1869, N920);
  xor KeyGate_0_24(KeyNOTWire_0[14], keyIn_0_24, KeyWire_0[24]);
  not KeyNOTGate_0_14(N1921, KeyNOTWire_0[14]);
  not NOT1_577 (KeyWire_0[25], N1869);
  xor KeyGate_0_25(KeyNOTWire_0[15], keyIn_0_25, KeyWire_0[25]);
  not KeyNOTGate_0_15(N1922, KeyNOTWire_0[15]);
not NOT1_578 (N1923, N1875);
nand NAND2_579 (N1924, N1714, N1895);
buf BUFF1_580 (N1927, N1858);
buf BUFF1_581 (N1930, N1858);
nand NAND2_582 (N1933, N1865, N1897);
nand NAND2_583 (N1936, N1882, N1911);
  not NOT1_584 (KeyWire_0[26], N1898);
  xor KeyGate_0_26(KeyNOTWire_0[16], keyIn_0_26, KeyWire_0[26]);
  not KeyNOTGate_0_16(N1937, KeyNOTWire_0[16]);
not NOT1_585 (N1938, N1902);
nand NAND2_586 (N1941, N679, N1920);
  nand NAND2_587 (KeyWire_0[27], N676, N1922);
  xor KeyGate_0_27(N1942, keyIn_0_27, KeyWire_0[27]);
buf BUFF1_588 (N1944, N1879);
not NOT1_589 (N1947, N1913);
buf BUFF1_590 (N1950, N1889);
buf BUFF1_591 (N1953, N1889);
buf BUFF1_592 (N1958, N1879);
nand NAND2_593 (N1961, N1896, N1924);
and AND2_594 (N1965, N1910, N601);
and AND2_595 (N1968, N602, N1912);
nand NAND2_596 (N1975, N1930, N917);
not NOT1_597 (N1976, N1930);
  nand NAND2_598 (KeyWire_0[28], N1927, N918);
  xor KeyGate_0_28(N1977, keyIn_0_28, KeyWire_0[28]);
  not NOT1_599 (KeyWire_0[29], N1927);
  xor KeyGate_0_29(KeyNOTWire_0[17], keyIn_0_29, KeyWire_0[29]);
  not KeyNOTGate_0_17(N1978, KeyNOTWire_0[17]);
nand NAND2_600 (N1979, N1919, N1941);
  nand NAND2_601 (KeyWire_0[30], N1921, N1942);
  xnor KeyGate_0_30(KeyNOTWire_0[18], keyIn_0_30, KeyWire_0[30]);
  not KeyNOTGate_0_18(N1980, KeyNOTWire_0[18]);
not NOT1_602 (N1985, N1933);
not NOT1_603 (N1987, N1936);
not NOT1_604 (N1999, N1944);
nand NAND2_605 (N2000, N1944, N1937);
not NOT1_606 (N2002, N1947);
nand NAND2_607 (N2003, N1947, N1499);
nand NAND2_608 (N2004, N1953, N1350);
not NOT1_609 (N2005, N1953);
  nand NAND2_610 (KeyWire_0[31], N1950, N1351);
  xnor KeyGate_0_31(KeyNOTWire_0[19], keyIn_0_31, KeyWire_0[31]);
  not KeyNOTGate_0_19(N2006, KeyNOTWire_0[19]);
  not NOT1_611 (KeyWire_0[32], N1950);
  xor KeyGate_0_32(KeyNOTWire_0[20], keyIn_0_32, KeyWire_0[32]);
  not KeyNOTGate_0_20(N2007, KeyNOTWire_0[20]);
nand NAND2_612 (N2008, N673, N1976);
  nand NAND2_613 (KeyWire_0[33], N670, N1978);
  xor KeyGate_0_33(KeyNOTWire_0[21], keyIn_0_33, KeyWire_0[33]);
  not KeyNOTGate_0_21(N2009, KeyNOTWire_0[21]);
not NOT1_614 (N2012, N1979);
not NOT1_615 (N2013, N1958);
nand NAND2_616 (N2014, N1958, N1923);
not NOT1_617 (N2015, N1961);
nand NAND2_618 (N2016, N1961, N1635);
not NOT1_619 (N2018, N1965);
not NOT1_620 (N2019, N1968);
nand NAND2_621 (N2020, N1898, N1999);
not NOT1_622 (N2021, N1987);
nand NAND2_623 (N2022, N1987, N1591);
nand NAND2_624 (N2023, N1440, N2002);
nand NAND2_625 (N2024, N1261, N2005);
  nand NAND2_626 (KeyWire_0[34], N1258, N2007);
  xor KeyGate_0_34(KeyNOTWire_0[22], keyIn_0_34, KeyWire_0[34]);
  not KeyNOTGate_0_22(N2025, KeyNOTWire_0[22]);
nand NAND2_627 (N2026, N1975, N2008);
  nand NAND2_628 (KeyWire_0[35], N1977, N2009);
  xor KeyGate_0_35(N2027, keyIn_0_35, KeyWire_0[35]);
  not NOT1_629 (KeyWire_0[36], N1980);
  xor KeyGate_0_36(KeyNOTWire_0[23], keyIn_0_36, KeyWire_0[36]);
  not KeyNOTGate_0_23(N2030, KeyNOTWire_0[23]);
buf BUFF1_630 (N2033, N1980);
nand NAND2_631 (N2036, N1875, N2013);
nand NAND2_632 (N2037, N1571, N2015);
nand NAND2_633 (N2038, N2020, N2000);
nand NAND2_634 (N2039, N1534, N2021);
nand NAND2_635 (N2040, N2023, N2003);
nand NAND2_636 (N2041, N2004, N2024);
  nand NAND2_637 (KeyWire_0[37], N2006, N2025);
  xor KeyGate_0_37(KeyNOTWire_0[24], keyIn_0_37, KeyWire_0[37]);
  not KeyNOTGate_0_24(N2042, KeyNOTWire_0[24]);
not NOT1_638 (N2047, N2026);
nand NAND2_639 (N2052, N2036, N2014);
nand NAND2_640 (N2055, N2037, N2016);
not NOT1_641 (N2060, N2038);
nand NAND2_642 (N2061, N2039, N2022);
nand NAND2_643 (N2062, N2040, N290);
not NOT1_644 (N2067, N2041);
  not NOT1_645 (KeyWire_0[38], N2027);
  xor KeyGate_0_38(N2068, keyIn_0_38, KeyWire_0[38]);
buf BUFF1_646 (N2071, N2027);
not NOT1_647 (N2076, N2052);
not NOT1_648 (N2077, N2055);
nand NAND2_649 (N2078, N2060, N290);
nand NAND2_650 (N2081, N2061, N290);
  not NOT1_651 (KeyWire_0[39], N2042);
  xor KeyGate_0_39(N2086, keyIn_0_39, KeyWire_0[39]);
buf BUFF1_652 (N2089, N2042);
  and AND2_653 (KeyWire_0[40], N2030, N2068);
  xor KeyGate_0_40(N2104, keyIn_0_40, KeyWire_0[40]);
  and AND2_654 (KeyWire_0[41], N2033, N2068);
  xor KeyGate_0_41(KeyNOTWire_0[25], keyIn_0_41, KeyWire_0[41]);
  not KeyNOTGate_0_25(N2119, KeyNOTWire_0[25]);
  and AND2_655 (KeyWire_0[42], N2030, N2071);
  xor KeyGate_0_42(KeyNOTWire_0[26], keyIn_0_42, KeyWire_0[42]);
  not KeyNOTGate_0_26(N2129, KeyNOTWire_0[26]);
and AND2_656 (N2143, N2033, N2071);
buf BUFF1_657 (N2148, N2062);
buf BUFF1_658 (N2151, N2062);
buf BUFF1_659 (N2196, N2078);
buf BUFF1_660 (N2199, N2078);
buf BUFF1_661 (N2202, N2081);
buf BUFF1_662 (N2205, N2081);
nand NAND2_663 (N2214, N2151, N915);
not NOT1_664 (N2215, N2151);
  nand NAND2_665 (KeyWire_0[43], N2148, N916);
  xor KeyGate_0_43(KeyNOTWire_0[27], keyIn_0_43, KeyWire_0[43]);
  not KeyNOTGate_0_27(N2216, KeyNOTWire_0[27]);
  not NOT1_666 (KeyWire_0[44], N2148);
  xor KeyGate_0_44(N2217, keyIn_0_44, KeyWire_0[44]);
nand NAND2_667 (N2222, N2199, N1348);
not NOT1_668 (N2223, N2199);
  nand NAND2_669 (KeyWire_0[45], N2196, N1349);
  xor KeyGate_0_45(KeyNOTWire_0[28], keyIn_0_45, KeyWire_0[45]);
  not KeyNOTGate_0_28(N2224, KeyNOTWire_0[28]);
  not NOT1_670 (KeyWire_0[46], N2196);
  xor KeyGate_0_46(N2225, keyIn_0_46, KeyWire_0[46]);
nand NAND2_671 (N2226, N2205, N913);
not NOT1_672 (N2227, N2205);
  nand NAND2_673 (KeyWire_0[47], N2202, N914);
  xnor KeyGate_0_47(N2228, keyIn_0_47, KeyWire_0[47]);
  not NOT1_674 (KeyWire_0[48], N2202);
  xor KeyGate_0_48(N2229, keyIn_0_48, KeyWire_0[48]);
nand NAND2_675 (N2230, N667, N2215);
  nand NAND2_676 (KeyWire_0[49], N664, N2217);
  xor KeyGate_0_49(N2231, keyIn_0_49, KeyWire_0[49]);
nand NAND2_677 (N2232, N1255, N2223);
  nand NAND2_678 (KeyWire_0[50], N1252, N2225);
  xor KeyGate_0_50(KeyNOTWire_0[29], keyIn_0_50, KeyWire_0[50]);
  not KeyNOTGate_0_29(N2233, KeyNOTWire_0[29]);
nand NAND2_679 (N2234, N661, N2227);
  nand NAND2_680 (KeyWire_0[51], N658, N2229);
  xnor KeyGate_0_51(KeyNOTWire_0[30], keyIn_0_51, KeyWire_0[51]);
  not KeyNOTGate_0_30(N2235, KeyNOTWire_0[30]);
nand NAND2_681 (N2236, N2214, N2230);
  nand NAND2_682 (KeyWire_0[52], N2216, N2231);
  xnor KeyGate_0_52(KeyNOTWire_0[31], keyIn_0_52, KeyWire_0[52]);
  not KeyNOTGate_0_31(N2237, KeyNOTWire_0[31]);
nand NAND2_683 (N2240, N2222, N2232);
  nand NAND2_684 (KeyWire_0[53], N2224, N2233);
  xnor KeyGate_0_53(N2241, keyIn_0_53, KeyWire_0[53]);
nand NAND2_685 (N2244, N2226, N2234);
  nand NAND2_686 (KeyWire_0[54], N2228, N2235);
  xor KeyGate_0_54(KeyNOTWire_0[32], keyIn_0_54, KeyWire_0[54]);
  not KeyNOTGate_0_32(N2245, KeyNOTWire_0[32]);
not NOT1_687 (N2250, N2236);
not NOT1_688 (N2253, N2240);
not NOT1_689 (N2256, N2244);
  not NOT1_690 (KeyWire_0[55], N2237);
  xor KeyGate_0_55(N2257, keyIn_0_55, KeyWire_0[55]);
buf BUFF1_691 (N2260, N2237);
  not NOT1_692 (KeyWire_0[56], N2241);
  xor KeyGate_0_56(KeyNOTWire_0[33], keyIn_0_56, KeyWire_0[56]);
  not KeyNOTGate_0_33(N2263, KeyNOTWire_0[33]);
and AND2_693 (N2266, N1164, N2241);
  not NOT1_694 (KeyWire_0[57], N2245);
  xor KeyGate_0_57(N2269, keyIn_0_57, KeyWire_0[57]);
and AND2_695 (N2272, N1168, N2245);
nand NAND8_696 (N2279, N2067, N2012, N2047, N2250, N899, N2256, N2253, N903);
buf BUFF1_697 (N2286, N2266);
buf BUFF1_698 (N2297, N2266);
buf BUFF1_699 (N2315, N2272);
buf BUFF1_700 (N2326, N2272);
  and AND2_701 (KeyWire_0[58], N2086, N2257);
  xnor KeyGate_0_58(N2340, keyIn_0_58, KeyWire_0[58]);
  and AND2_702 (KeyWire_0[59], N2089, N2257);
  xnor KeyGate_0_59(N2353, keyIn_0_59, KeyWire_0[59]);
  and AND2_703 (KeyWire_0[60], N2086, N2260);
  xor KeyGate_0_60(KeyNOTWire_0[34], keyIn_0_60, KeyWire_0[60]);
  not KeyNOTGate_0_34(N2361, KeyNOTWire_0[34]);
  and AND2_704 (KeyWire_0[61], N2089, N2260);
  xor KeyGate_0_61(KeyNOTWire_0[35], keyIn_0_61, KeyWire_0[61]);
  not KeyNOTGate_0_35(N2375, KeyNOTWire_0[35]);
and AND4_705 (N2384, N338, N2279, N313, N313);
and AND2_706 (N2385, N1163, N2263);
  and AND2_707 (KeyWire_0[62], N1164, N2263);
  xnor KeyGate_0_62(N2386, keyIn_0_62, KeyWire_0[62]);
and AND2_708 (N2426, N1167, N2269);
  and AND2_709 (KeyWire_0[63], N1168, N2269);
  xor KeyGate_0_63(N2427, keyIn_0_63, KeyWire_0[63]);
  nand NAND5_710 (KeyWire_0[64], N2286, N2315, N2361, N2104, N1171);
  xnor KeyGate_0_64(N2537, keyIn_0_64, KeyWire_0[64]);
  nand NAND5_711 (KeyWire_0[65], N2286, N2315, N2340, N2129, N1171);
  xor KeyGate_0_65(KeyNOTWire_0[36], keyIn_0_65, KeyWire_0[65]);
  not KeyNOTGate_0_36(N2540, KeyNOTWire_0[36]);
  nand NAND5_712 (KeyWire_0[66], N2286, N2315, N2340, N2119, N1171);
  xnor KeyGate_0_66(KeyNOTWire_0[37], keyIn_0_66, KeyWire_0[66]);
  not KeyNOTGate_0_37(N2543, KeyNOTWire_0[37]);
  nand NAND5_713 (KeyWire_0[67], N2286, N2315, N2353, N2104, N1171);
  xnor KeyGate_0_67(KeyNOTWire_0[38], keyIn_0_67, KeyWire_0[67]);
  not KeyNOTGate_0_38(N2546, KeyNOTWire_0[38]);
  nand NAND5_714 (KeyWire_0[68], N2297, N2315, N2375, N2119, N1188);
  xor KeyGate_0_68(N2549, keyIn_0_68, KeyWire_0[68]);
  nand NAND5_715 (KeyWire_0[69], N2297, N2326, N2361, N2143, N1188);
  xnor KeyGate_0_69(N2552, keyIn_0_69, KeyWire_0[69]);
  nand NAND5_716 (KeyWire_0[70], N2297, N2326, N2375, N2129, N1188);
  xor KeyGate_0_70(KeyNOTWire_0[39], keyIn_0_70, KeyWire_0[70]);
  not KeyNOTGate_0_39(N2555, KeyNOTWire_0[39]);
and AND5_717 (N2558, N2286, N2315, N2361, N2104, N1171);
and AND5_718 (N2561, N2286, N2315, N2340, N2129, N1171);
and AND5_719 (N2564, N2286, N2315, N2340, N2119, N1171);
and AND5_720 (N2567, N2286, N2315, N2353, N2104, N1171);
and AND5_721 (N2570, N2297, N2315, N2375, N2119, N1188);
and AND5_722 (N2573, N2297, N2326, N2361, N2143, N1188);
and AND5_723 (N2576, N2297, N2326, N2375, N2129, N1188);
  nand NAND5_724 (KeyWire_0[71], N2286, N2427, N2361, N2129, N1171);
  xor KeyGate_0_71(KeyNOTWire_0[40], keyIn_0_71, KeyWire_0[71]);
  not KeyNOTGate_0_40(N2594, KeyNOTWire_0[40]);
  nand NAND5_725 (KeyWire_0[72], N2297, N2427, N2361, N2119, N1171);
  xnor KeyGate_0_72(N2597, keyIn_0_72, KeyWire_0[72]);
  nand NAND5_726 (KeyWire_0[73], N2297, N2427, N2375, N2104, N1171);
  xnor KeyGate_0_73(KeyNOTWire_0[41], keyIn_0_73, KeyWire_0[73]);
  not KeyNOTGate_0_41(N2600, KeyNOTWire_0[41]);
  nand NAND5_727 (KeyWire_0[74], N2297, N2427, N2340, N2143, N1171);
  xnor KeyGate_0_74(KeyNOTWire_0[42], keyIn_0_74, KeyWire_0[74]);
  not KeyNOTGate_0_42(N2603, KeyNOTWire_0[42]);
  nand NAND5_728 (KeyWire_0[75], N2297, N2427, N2353, N2129, N1188);
  xor KeyGate_0_75(KeyNOTWire_0[43], keyIn_0_75, KeyWire_0[75]);
  not KeyNOTGate_0_43(N2606, KeyNOTWire_0[43]);
  nand NAND5_729 (KeyWire_0[76], N2386, N2326, N2361, N2129, N1188);
  xor KeyGate_0_76(N2611, keyIn_0_76, KeyWire_0[76]);
  nand NAND5_730 (KeyWire_0[77], N2386, N2326, N2361, N2119, N1188);
  xnor KeyGate_0_77(KeyNOTWire_0[44], keyIn_0_77, KeyWire_0[77]);
  not KeyNOTGate_0_44(N2614, KeyNOTWire_0[44]);
  nand NAND5_731 (KeyWire_0[78], N2386, N2326, N2375, N2104, N1188);
  xnor KeyGate_0_78(N2617, keyIn_0_78, KeyWire_0[78]);
  nand NAND5_732 (KeyWire_0[79], N2386, N2326, N2353, N2129, N1188);
  xor KeyGate_0_79(N2620, keyIn_0_79, KeyWire_0[79]);
nand NAND5_733 (N2627, N2297, N2427, N2340, N2104, N926);
nand NAND5_734 (N2628, N2386, N2326, N2340, N2104, N926);
nand NAND5_735 (N2629, N2386, N2427, N2361, N2104, N926);
nand NAND5_736 (N2630, N2386, N2427, N2340, N2129, N926);
nand NAND5_737 (N2631, N2386, N2427, N2340, N2119, N926);
nand NAND5_738 (N2632, N2386, N2427, N2353, N2104, N926);
nand NAND5_739 (N2633, N2386, N2426, N2340, N2104, N926);
nand NAND5_740 (N2634, N2385, N2427, N2340, N2104, N926);
and AND5_741 (N2639, N2286, N2427, N2361, N2129, N1171);
and AND5_742 (N2642, N2297, N2427, N2361, N2119, N1171);
and AND5_743 (N2645, N2297, N2427, N2375, N2104, N1171);
and AND5_744 (N2648, N2297, N2427, N2340, N2143, N1171);
and AND5_745 (N2651, N2297, N2427, N2353, N2129, N1188);
and AND5_746 (N2655, N2386, N2326, N2361, N2129, N1188);
and AND5_747 (N2658, N2386, N2326, N2361, N2119, N1188);
and AND5_748 (N2661, N2386, N2326, N2375, N2104, N1188);
and AND5_749 (N2664, N2386, N2326, N2353, N2129, N1188);
nand NAND2_750 (N2669, N2558, N534);
not NOT1_751 (N2670, N2558);
nand NAND2_752 (N2671, N2561, N535);
not NOT1_753 (N2672, N2561);
nand NAND2_754 (N2673, N2564, N536);
not NOT1_755 (N2674, N2564);
nand NAND2_756 (N2675, N2567, N537);
not NOT1_757 (N2676, N2567);
nand NAND2_758 (N2682, N2570, N543);
not NOT1_759 (N2683, N2570);
nand NAND2_760 (N2688, N2573, N548);
not NOT1_761 (N2689, N2573);
nand NAND2_762 (N2690, N2576, N549);
not NOT1_763 (N2691, N2576);
and AND8_764 (N2710, N2627, N2628, N2629, N2630, N2631, N2632, N2633, N2634);
nand NAND2_765 (N2720, N343, N2670);
nand NAND2_766 (N2721, N346, N2672);
nand NAND2_767 (N2722, N349, N2674);
nand NAND2_768 (N2723, N352, N2676);
nand NAND2_769 (N2724, N2639, N538);
not NOT1_770 (N2725, N2639);
nand NAND2_771 (N2726, N2642, N539);
not NOT1_772 (N2727, N2642);
  nand NAND2_773 (KeyWire_0[80], N2645, N540);
  xor KeyGate_0_80(KeyNOTWire_0[45], keyIn_0_80, KeyWire_0[80]);
  not KeyNOTGate_0_45(N2728, KeyNOTWire_0[45]);
not NOT1_774 (N2729, N2645);
nand NAND2_775 (N2730, N2648, N541);
not NOT1_776 (N2731, N2648);
nand NAND2_777 (N2732, N2651, N542);
not NOT1_778 (N2733, N2651);
nand NAND2_779 (N2734, N370, N2683);
nand NAND2_780 (N2735, N2655, N544);
not NOT1_781 (N2736, N2655);
nand NAND2_782 (N2737, N2658, N545);
not NOT1_783 (N2738, N2658);
nand NAND2_784 (N2739, N2661, N546);
not NOT1_785 (N2740, N2661);
nand NAND2_786 (N2741, N2664, N547);
not NOT1_787 (N2742, N2664);
nand NAND2_788 (N2743, N385, N2689);
nand NAND2_789 (N2744, N388, N2691);
nand NAND8_790 (N2745, N2537, N2540, N2543, N2546, N2594, N2597, N2600, N2603);
nand NAND8_791 (N2746, N2606, N2549, N2611, N2614, N2617, N2620, N2552, N2555);
  and AND8_792 (KeyWire_0[81], N2537, N2540, N2543, N2546, N2594, N2597, N2600, N2603);
  xor KeyGate_0_81(KeyNOTWire_0[46], keyIn_0_81, KeyWire_0[81]);
  not KeyNOTGate_0_46(N2747, KeyNOTWire_0[46]);
  and AND8_793 (KeyWire_0[82], N2606, N2549, N2611, N2614, N2617, N2620, N2552, N2555);
  xnor KeyGate_0_82(KeyNOTWire_0[47], keyIn_0_82, KeyWire_0[82]);
  not KeyNOTGate_0_47(N2750, KeyNOTWire_0[47]);
nand NAND2_794 (N2753, N2669, N2720);
nand NAND2_795 (N2754, N2671, N2721);
nand NAND2_796 (N2755, N2673, N2722);
nand NAND2_797 (N2756, N2675, N2723);
nand NAND2_798 (N2757, N355, N2725);
nand NAND2_799 (N2758, N358, N2727);
nand NAND2_800 (N2759, N361, N2729);
nand NAND2_801 (N2760, N364, N2731);
nand NAND2_802 (N2761, N367, N2733);
nand NAND2_803 (N2762, N2682, N2734);
nand NAND2_804 (N2763, N373, N2736);
nand NAND2_805 (N2764, N376, N2738);
nand NAND2_806 (N2765, N379, N2740);
nand NAND2_807 (N2766, N382, N2742);
nand NAND2_808 (N2767, N2688, N2743);
nand NAND2_809 (N2768, N2690, N2744);
and AND2_810 (N2773, N2745, N275);
and AND2_811 (N2776, N2746, N276);
nand NAND2_812 (N2779, N2724, N2757);
nand NAND2_813 (N2780, N2726, N2758);
nand NAND2_814 (N2781, N2728, N2759);
nand NAND2_815 (N2782, N2730, N2760);
nand NAND2_816 (N2783, N2732, N2761);
nand NAND2_817 (N2784, N2735, N2763);
nand NAND2_818 (N2785, N2737, N2764);
nand NAND2_819 (N2786, N2739, N2765);
nand NAND2_820 (N2787, N2741, N2766);
  and AND3_821 (KeyWire_0[83], N2747, N2750, N2710);
  xnor KeyGate_0_83(KeyNOTWire_0[48], keyIn_0_83, KeyWire_0[83]);
  not KeyNOTGate_0_48(N2788, KeyNOTWire_0[48]);
  nand NAND2_822 (KeyWire_0[84], N2747, N2750);
  xor KeyGate_0_84(N2789, keyIn_0_84, KeyWire_0[84]);
  and AND4_823 (KeyWire_0[85], N338, N2279, N99, N2788);
  xor KeyGate_0_85(N2800, keyIn_0_85, KeyWire_0[85]);
nand NAND2_824 (N2807, N2773, N2018);
not NOT1_825 (N2808, N2773);
nand NAND2_826 (N2809, N2776, N2019);
not NOT1_827 (N2810, N2776);
  nor NOR2_828 (KeyWire_0[86], N2384, N2800);
  xnor KeyGate_0_86(KeyNOTWire_0[49], keyIn_0_86, KeyWire_0[86]);
  not KeyNOTGate_0_49(N2811, KeyNOTWire_0[49]);
  and AND3_829 (KeyWire_0[87], N897, N283, N2789);
  xnor KeyGate_0_87(KeyNOTWire_0[50], keyIn_0_87, KeyWire_0[87]);
  not KeyNOTGate_0_50(N2812, KeyNOTWire_0[50]);
  and AND3_830 (KeyWire_0[88], N76, N283, N2789);
  xnor KeyGate_0_88(N2815, keyIn_0_88, KeyWire_0[88]);
  and AND3_831 (KeyWire_0[89], N82, N283, N2789);
  xnor KeyGate_0_89(N2818, keyIn_0_89, KeyWire_0[89]);
  and AND3_832 (KeyWire_0[90], N85, N283, N2789);
  xor KeyGate_0_90(KeyNOTWire_0[51], keyIn_0_90, KeyWire_0[90]);
  not KeyNOTGate_0_51(N2821, KeyNOTWire_0[51]);
  and AND3_833 (KeyWire_0[91], N898, N283, N2789);
  xnor KeyGate_0_91(KeyNOTWire_0[52], keyIn_0_91, KeyWire_0[91]);
  not KeyNOTGate_0_52(N2824, KeyNOTWire_0[52]);
nand NAND2_834 (N2827, N1965, N2808);
nand NAND2_835 (N2828, N1968, N2810);
  and AND3_836 (KeyWire_0[92], N79, N283, N2789);
  xnor KeyGate_0_92(KeyNOTWire_0[53], keyIn_0_92, KeyWire_0[92]);
  not KeyNOTGate_0_53(N2829, KeyNOTWire_0[53]);
nand NAND2_837 (N2843, N2807, N2827);
  nand NAND2_838 (KeyWire_0[93], N2809, N2828);
  xnor KeyGate_0_93(N2846, keyIn_0_93, KeyWire_0[93]);
  nand NAND2_839 (KeyWire_0[94], N2812, N2076);
  xor KeyGate_0_94(KeyNOTWire_0[54], keyIn_0_94, KeyWire_0[94]);
  not KeyNOTGate_0_54(N2850, KeyNOTWire_0[54]);
  nand NAND2_840 (KeyWire_0[95], N2815, N2077);
  xnor KeyGate_0_95(KeyNOTWire_0[55], keyIn_0_95, KeyWire_0[95]);
  not KeyNOTGate_0_55(N2851, KeyNOTWire_0[55]);
  nand NAND2_841 (KeyWire_0[96], N2818, N1915);
  xnor KeyGate_0_96(N2852, keyIn_0_96, KeyWire_0[96]);
  nand NAND2_842 (KeyWire_0[97], N2821, N1857);
  xor KeyGate_0_97(KeyNOTWire_0[56], keyIn_0_97, KeyWire_0[97]);
  not KeyNOTGate_0_56(N2853, KeyNOTWire_0[56]);
  nand NAND2_843 (KeyWire_0[98], N2824, N1938);
  xnor KeyGate_0_98(N2854, keyIn_0_98, KeyWire_0[98]);
  not NOT1_844 (KeyWire_0[99], N2812);
  xnor KeyGate_0_99(KeyNOTWire_0[57], keyIn_0_99, KeyWire_0[99]);
  not KeyNOTGate_0_57(N2857, KeyNOTWire_0[57]);
  not NOT1_845 (KeyWire_0[100], N2815);
  xnor KeyGate_0_100(N2858, keyIn_0_100, KeyWire_0[100]);
  not NOT1_846 (KeyWire_0[101], N2818);
  xor KeyGate_0_101(KeyNOTWire_0[58], keyIn_0_101, KeyWire_0[101]);
  not KeyNOTGate_0_58(N2859, KeyNOTWire_0[58]);
  not NOT1_847 (KeyWire_0[102], N2821);
  xor KeyGate_0_102(KeyNOTWire_0[59], keyIn_0_102, KeyWire_0[102]);
  not KeyNOTGate_0_59(N2860, KeyNOTWire_0[59]);
  not NOT1_848 (KeyWire_0[103], N2824);
  xnor KeyGate_0_103(KeyNOTWire_0[60], keyIn_0_103, KeyWire_0[103]);
  not KeyNOTGate_0_60(N2861, KeyNOTWire_0[60]);
  not NOT1_849 (KeyWire_0[104], N2829);
  xor KeyGate_0_104(N2862, keyIn_0_104, KeyWire_0[104]);
  nand NAND2_850 (KeyWire_0[105], N2829, N1985);
  xor KeyGate_0_105(N2863, keyIn_0_105, KeyWire_0[105]);
  nand NAND2_851 (KeyWire_0[106], N2052, N2857);
  xnor KeyGate_0_106(N2866, keyIn_0_106, KeyWire_0[106]);
  nand NAND2_852 (KeyWire_0[107], N2055, N2858);
  xnor KeyGate_0_107(KeyNOTWire_0[61], keyIn_0_107, KeyWire_0[107]);
  not KeyNOTGate_0_61(N2867, KeyNOTWire_0[61]);
  nand NAND2_853 (KeyWire_0[108], N1866, N2859);
  xnor KeyGate_0_108(N2868, keyIn_0_108, KeyWire_0[108]);
  nand NAND2_854 (KeyWire_0[109], N1818, N2860);
  xor KeyGate_0_109(KeyNOTWire_0[62], keyIn_0_109, KeyWire_0[109]);
  not KeyNOTGate_0_62(N2869, KeyNOTWire_0[62]);
  nand NAND2_855 (KeyWire_0[110], N1902, N2861);
  xnor KeyGate_0_110(KeyNOTWire_0[63], keyIn_0_110, KeyWire_0[110]);
  not KeyNOTGate_0_63(N2870, KeyNOTWire_0[63]);
nand NAND2_856 (N2871, N2843, N886);
not NOT1_857 (N2872, N2843);
nand NAND2_858 (N2873, N2846, N887);
not NOT1_859 (N2874, N2846);
  nand NAND2_860 (KeyWire_0[111], N1933, N2862);
  xnor KeyGate_0_111(N2875, keyIn_0_111, KeyWire_0[111]);
  nand NAND2_861 (KeyWire_0[112], N2866, N2850);
  xnor KeyGate_0_112(N2876, keyIn_0_112, KeyWire_0[112]);
  nand NAND2_862 (KeyWire_0[113], N2867, N2851);
  xnor KeyGate_0_113(N2877, keyIn_0_113, KeyWire_0[113]);
  nand NAND2_863 (KeyWire_0[114], N2868, N2852);
  xnor KeyGate_0_114(N2878, keyIn_0_114, KeyWire_0[114]);
  nand NAND2_864 (KeyWire_0[115], N2869, N2853);
  xnor KeyGate_0_115(KeyNOTWire_0[64], keyIn_0_115, KeyWire_0[115]);
  not KeyNOTGate_0_64(N2879, KeyNOTWire_0[64]);
  nand NAND2_865 (KeyWire_0[116], N2870, N2854);
  xor KeyGate_0_116(N2880, keyIn_0_116, KeyWire_0[116]);
nand NAND2_866 (N2881, N682, N2872);
nand NAND2_867 (N2882, N685, N2874);
  nand NAND2_868 (KeyWire_0[117], N2875, N2863);
  xnor KeyGate_0_117(KeyNOTWire_0[65], keyIn_0_117, KeyWire_0[117]);
  not KeyNOTGate_0_65(N2883, KeyNOTWire_0[65]);
  and AND2_869 (KeyWire_0[118], N2876, N550);
  xnor KeyGate_0_118(KeyNOTWire_0[66], keyIn_0_118, KeyWire_0[118]);
  not KeyNOTGate_0_66(N2886, KeyNOTWire_0[66]);
  and AND2_870 (KeyWire_0[119], N551, N2877);
  xnor KeyGate_0_119(KeyNOTWire_0[67], keyIn_0_119, KeyWire_0[119]);
  not KeyNOTGate_0_67(N2887, KeyNOTWire_0[67]);
  and AND2_871 (KeyWire_0[120], N553, N2878);
  xor KeyGate_0_120(KeyNOTWire_0[68], keyIn_0_120, KeyWire_0[120]);
  not KeyNOTGate_0_68(N2888, KeyNOTWire_0[68]);
  and AND2_872 (KeyWire_0[121], N2879, N554);
  xor KeyGate_0_121(N2889, keyIn_0_121, KeyWire_0[121]);
  and AND2_873 (KeyWire_0[122], N555, N2880);
  xor KeyGate_0_122(KeyNOTWire_0[69], keyIn_0_122, KeyWire_0[122]);
  not KeyNOTGate_0_69(N2890, KeyNOTWire_0[69]);
nand NAND2_874 (N2891, N2871, N2881);
nand NAND2_875 (N2892, N2873, N2882);
  nand NAND2_876 (KeyWire_0[123], N2883, N1461);
  xor KeyGate_0_123(KeyNOTWire_0[70], keyIn_0_123, KeyWire_0[123]);
  not KeyNOTGate_0_70(N2895, KeyNOTWire_0[70]);
  not NOT1_877 (KeyWire_0[124], N2883);
  xnor KeyGate_0_124(N2896, keyIn_0_124, KeyWire_0[124]);
  nand NAND2_878 (KeyWire_0[125], N1383, N2896);
  xnor KeyGate_0_125(N2897, keyIn_0_125, KeyWire_0[125]);
  nand NAND2_879 (KeyWire_0[126], N2895, N2897);
  xnor KeyGate_0_126(KeyNOTWire_0[71], keyIn_0_126, KeyWire_0[126]);
  not KeyNOTGate_0_71(N2898, KeyNOTWire_0[71]);
  and AND2_880 (KeyWire_0[127], N2898, N552);
  xnor KeyGate_0_127(N2899, keyIn_0_127, KeyWire_0[127]);

endmodule
