// Verilog File 
module top (G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,
G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,
G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,
G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat,G223gat,G329gat,G370gat,
G421gat,G430gat,G431gat,G432gat,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,
keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,
keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,
keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,keyinput35,
keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,keyinput45,
keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,keyinput55,
keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,keyinput65,
keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,keyinput75,
keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,keyinput85,
keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,keyinput95,
keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,keyinput105,
keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,keyinput115,
keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,keyinput125,
keyinput126,keyinput127,keyinput128,keyinput129,keyinput130,keyinput131,keyinput132,keyinput133,keyinput134,keyinput135,
keyinput136,keyinput137,keyinput138,keyinput139,keyinput140,keyinput141,keyinput142,keyinput143,keyinput144,keyinput145,
keyinput146,keyinput147,keyinput148,keyinput149,keyinput150,keyinput151,keyinput152,keyinput153,keyinput154,keyinput155,
keyinput156,keyinput157,keyinput158,keyinput159,keyinput160,keyinput161,keyinput162,keyinput163,keyinput164,keyinput165,
keyinput166,keyinput167,keyinput168,keyinput169,keyinput170,keyinput171,keyinput172,keyinput173,keyinput174,keyinput175,
keyinput176,keyinput177,keyinput178,keyinput179,keyinput180,keyinput181,keyinput182,keyinput183,keyinput184,keyinput185,
keyinput186,keyinput187,keyinput188,keyinput189,keyinput190,keyinput191,keyinput192,keyinput193,keyinput194,keyinput195,
keyinput196,keyinput197,keyinput198,keyinput199);

input G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,
G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,
G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,
G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat,keyinput0,keyinput1,keyinput2,
keyinput3,keyinput4,keyinput5,keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,
keyinput13,keyinput14,keyinput15,keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,
keyinput23,keyinput24,keyinput25,keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,
keyinput33,keyinput34,keyinput35,keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,
keyinput43,keyinput44,keyinput45,keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,
keyinput53,keyinput54,keyinput55,keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,
keyinput63,keyinput64,keyinput65,keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,
keyinput73,keyinput74,keyinput75,keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,
keyinput83,keyinput84,keyinput85,keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,
keyinput93,keyinput94,keyinput95,keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,
keyinput103,keyinput104,keyinput105,keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,
keyinput113,keyinput114,keyinput115,keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,
keyinput123,keyinput124,keyinput125,keyinput126,keyinput127,keyinput128,keyinput129,keyinput130,keyinput131,keyinput132,
keyinput133,keyinput134,keyinput135,keyinput136,keyinput137,keyinput138,keyinput139,keyinput140,keyinput141,keyinput142,
keyinput143,keyinput144,keyinput145,keyinput146,keyinput147,keyinput148,keyinput149,keyinput150,keyinput151,keyinput152,
keyinput153,keyinput154,keyinput155,keyinput156,keyinput157,keyinput158,keyinput159,keyinput160,keyinput161,keyinput162,
keyinput163,keyinput164,keyinput165,keyinput166,keyinput167,keyinput168,keyinput169,keyinput170,keyinput171,keyinput172,
keyinput173,keyinput174,keyinput175,keyinput176,keyinput177,keyinput178,keyinput179,keyinput180,keyinput181,keyinput182,
keyinput183,keyinput184,keyinput185,keyinput186,keyinput187,keyinput188,keyinput189,keyinput190,keyinput191,keyinput192,
keyinput193,keyinput194,keyinput195,keyinput196,keyinput197,keyinput198,keyinput199;

output G223gat,G329gat,G370gat,G421gat,G430gat,G431gat,G432gat;

wire G118gat,G119gat,G122gat,G123gat,G126gat,G127gat,G130gat,G131gat,G134gat,
G135gat,G138gat,G139gat,G142gat,G143gat,G146gat,G147gat,G150gat,G151gat,G154gat,
G157gat,G158gat,G159gat,G162gat,G165gat,G168gat,G171gat,G174gat,G177gat,G180gat,
G183gat,G184gat,G185gat,G186gat,G187gat,G188gat,G189gat,G190gat,G191gat,G192gat,
G193gat,G194gat,G195gat,G196gat,G197gat,G198gat,G199gat,G203gat,G213gat,G224gat,
G227gat,G230gat,G233gat,G236gat,G239gat,G242gat,G243gat,G246gat,G247gat,G250gat,
G251gat,G254gat,G255gat,G256gat,G257gat,G258gat,G259gat,G260gat,G263gat,G264gat,
G267gat,G270gat,G273gat,G276gat,G279gat,G282gat,G285gat,G288gat,G289gat,G290gat,
G291gat,G292gat,G293gat,G294gat,G295gat,G296gat,G300gat,G301gat,G302gat,G303gat,
G304gat,G305gat,G306gat,G307gat,G308gat,G309gat,G319gat,G330gat,G331gat,G332gat,
G333gat,G334gat,G335gat,G336gat,G337gat,G338gat,G339gat,G340gat,G341gat,G342gat,
G343gat,G344gat,G345gat,G346gat,G347gat,G348gat,G349gat,G350gat,G351gat,G352gat,
G353gat,G354gat,G355gat,G356gat,G357gat,G360gat,G371gat,G372gat,G373gat,G374gat,
G375gat,G376gat,G377gat,G378gat,G379gat,G380gat,G381gat,G386gat,G393gat,G399gat,
G404gat,G407gat,G411gat,G414gat,G415gat,G416gat,G417gat,G418gat,G419gat,G420gat,
G422gat,G425gat,G428gat,G429gat,muxed0,muxed1,muxed2,muxed3,muxed4,muxed5,
muxed6,muxed7,muxed8,muxed9,muxed10,muxed11,muxed12,muxed13,muxed14,muxed15,
muxed16,muxed17,muxed18,muxed19,muxed20,muxed21,muxed22,muxed23,muxed24,muxed25,
muxed26,muxed27,muxed28,muxed29,muxed30,muxed31,muxed32,muxed33,muxed34,muxed35,
muxed36,muxed37,muxed38,muxed39,muxed40,muxed41,muxed42,muxed43,muxed44,muxed45,
muxed46,muxed47,muxed48,muxed49,muxed50,muxed51,muxed52,muxed53,muxed54,muxed55,
muxed56,muxed57,muxed58,muxed59,muxed60,muxed61,muxed62,muxed63,muxed64,muxed65,
muxed66,muxed67,muxed68,muxed69,muxed70,muxed71,muxed72,muxed73,muxed74,muxed75,
muxed76,muxed77,muxed78,muxed79,muxed80,muxed81,muxed82,muxed83,muxed84,muxed85,
muxed86,muxed87,muxed88,muxed89,muxed90,muxed91,muxed92,muxed93,muxed94,muxed95,
muxed96,muxed97,muxed98,muxed99,muxed100,muxed101,muxed102,muxed103,muxed104,muxed105,
muxed106,muxed107,muxed108,muxed109,muxed110,muxed111,muxed112,muxed113,muxed114,muxed115,
muxed116,muxed117,muxed118,muxed119,muxed120,muxed121,muxed122,muxed123,muxed124,muxed125,
muxed126,muxed127,muxed128,muxed129,muxed130,muxed131,muxed132,muxed133,muxed134,muxed135,
muxed136,muxed137,muxed138,muxed139,muxed140,muxed141,muxed142,muxed143,muxed144,muxed145,
muxed146,muxed147,muxed148,muxed149,muxed150,muxed151,muxed152,muxed153,muxed154,muxed155,
muxed156,muxed157,muxed158,muxed159,muxed160,muxed161,muxed162,muxed163,muxed164,muxed165,
muxed166,muxed167,muxed168,muxed169,muxed170,muxed171,muxed172,muxed173,muxed174,muxed175,
muxed176,muxed177,muxed178,muxed179,muxed180,muxed181,muxed182,muxed183,muxed184,muxed185,
muxed186,muxed187,muxed188,muxed189,muxed190,muxed191,muxed192,muxed193,muxed194,muxed195,
muxed196,muxed197,muxed198,muxed199;
not gate_0(G118gat,G1gat);
not gate_1(G119gat,G4gat);
not gate_2(G122gat,G11gat);
not gate_3(G123gat,G17gat);
not gate_4(G126gat,G24gat);
not gate_5(G127gat,G30gat);
not gate_6(G130gat,G37gat);
not gate_7(G131gat,muxed189);
not gate_8(G134gat,G50gat);
not gate_9(G135gat,G56gat);
not gate_10(G138gat,G63gat);
not gate_11(G139gat,G69gat);
not gate_12(G142gat,muxed14);
not gate_13(G143gat,G82gat);
not gate_14(G146gat,G89gat);
not gate_15(G147gat,G95gat);
not gate_16(G150gat,muxed186);
not gate_17(G151gat,G108gat);
nand gate_18(G154gat,G118gat,G4gat);
nor gate_19(G157gat,muxed66,muxed27);
nor gate_20(G158gat,G14gat,muxed27);
nand gate_21(G159gat,muxed158,G17gat);
nand gate_22(G162gat,muxed164,G30gat);
nand gate_23(G165gat,G130gat,muxed189);
nand gate_24(G168gat,G134gat,G56gat);
nand gate_25(G171gat,G138gat,G69gat);
nand gate_26(G174gat,muxed36,G82gat);
nand gate_27(G177gat,muxed3,G95gat);
nand gate_28(G180gat,muxed122,G108gat);
nor gate_29(G183gat,G21gat,G123gat);
nor gate_30(G184gat,G27gat,G123gat);
nor gate_31(G185gat,G34gat,muxed32);
nor gate_32(G186gat,G40gat,muxed32);
nor gate_33(G187gat,G47gat,muxed39);
nor gate_34(G188gat,G53gat,muxed39);
nor gate_35(G189gat,G60gat,muxed109);
nor gate_36(G190gat,G66gat,muxed109);
nor gate_37(G191gat,G73gat,G139gat);
nor gate_38(G192gat,G79gat,G139gat);
nor gate_39(G193gat,G86gat,G143gat);
nor gate_40(G194gat,G92gat,G143gat);
nor gate_41(G195gat,G99gat,G147gat);
nor gate_42(G196gat,G105gat,G147gat);
nor gate_43(G197gat,G112gat,G151gat);
nor gate_44(G198gat,G115gat,G151gat);
and gate_45(G199gat,G154gat,muxed97,muxed175,G165gat,G168gat,G171gat,muxed33,G177gat,muxed63);
not gate_46(G203gat,G199gat);
not gate_47(G213gat,G199gat);
not gate_48(G223gat,G199gat);
xor gate_49(G224gat,G203gat,G154gat);
xor gate_50(G227gat,G203gat,muxed97);
xor gate_51(G230gat,G203gat,muxed175);
xor gate_52(G233gat,G203gat,G165gat);
xor gate_53(G236gat,G203gat,G168gat);
xor gate_54(G239gat,G203gat,G171gat);
nand gate_55(G242gat,G1gat,muxed88);
xor gate_56(G243gat,G203gat,muxed33);
nand gate_57(G246gat,muxed88,G11gat);
xor gate_58(G247gat,G203gat,G177gat);
nand gate_59(G250gat,muxed88,G24gat);
xor gate_60(G251gat,G203gat,muxed63);
nand gate_61(G254gat,muxed88,G37gat);
nand gate_62(G255gat,muxed88,G50gat);
nand gate_63(G256gat,muxed88,G63gat);
nand gate_64(G257gat,muxed88,muxed14);
nand gate_65(G258gat,muxed88,G89gat);
nand gate_66(G259gat,muxed88,muxed186);
nand gate_67(G260gat,G224gat,muxed75);
nand gate_68(G263gat,G224gat,muxed194);
nand gate_69(G264gat,muxed0,G183gat);
nand gate_70(G267gat,muxed170,G185gat);
nand gate_71(G270gat,muxed114,G187gat);
nand gate_72(G273gat,muxed35,G189gat);
nand gate_73(G276gat,muxed188,G191gat);
nand gate_74(G279gat,muxed30,muxed180);
nand gate_75(G282gat,G247gat,G195gat);
nand gate_76(G285gat,muxed125,muxed147);
nand gate_77(G288gat,muxed0,muxed5);
nand gate_78(G289gat,muxed170,G186gat);
nand gate_79(G290gat,muxed114,muxed38);
nand gate_80(G291gat,muxed35,muxed183);
nand gate_81(G292gat,muxed188,G192gat);
nand gate_82(G293gat,muxed30,G194gat);
nand gate_83(G294gat,G247gat,G196gat);
nand gate_84(G295gat,muxed125,G198gat);
and gate_85(G296gat,muxed113,G264gat,G267gat,G270gat,G273gat,muxed11,G279gat,muxed23,muxed137);
not gate_86(G300gat,muxed192);
not gate_87(G301gat,muxed12);
not gate_88(G302gat,muxed50);
not gate_89(G303gat,muxed19);
not gate_90(G304gat,muxed178);
not gate_91(G305gat,muxed199);
not gate_92(G306gat,muxed22);
not gate_93(G307gat,muxed138);
not gate_94(G308gat,muxed100);
not gate_95(G309gat,muxed124);
not gate_96(G319gat,muxed124);
not gate_97(G329gat,muxed124);
xor gate_98(G330gat,muxed151,muxed113);
xor gate_99(G331gat,muxed151,G264gat);
xor gate_100(G332gat,muxed151,G267gat);
xor gate_101(G333gat,muxed151,G270gat);
nand gate_102(G334gat,muxed66,muxed123);
xor gate_103(G335gat,muxed151,G273gat);
nand gate_104(G336gat,muxed123,G21gat);
xor gate_105(G337gat,muxed151,muxed11);
nand gate_106(G338gat,muxed123,G34gat);
xor gate_107(G339gat,muxed151,G279gat);
nand gate_108(G340gat,muxed123,G47gat);
xor gate_109(G341gat,muxed151,muxed23);
nand gate_110(G342gat,muxed123,G60gat);
xor gate_111(G343gat,muxed151,muxed137);
nand gate_112(G344gat,muxed123,G73gat);
nand gate_113(G345gat,muxed123,G86gat);
nand gate_114(G346gat,muxed123,G99gat);
nand gate_115(G347gat,muxed123,G112gat);
nand gate_116(G348gat,muxed83,muxed191);
nand gate_117(G349gat,muxed21,muxed10);
nand gate_118(G350gat,G332gat,muxed70);
nand gate_119(G351gat,G333gat,G303gat);
nand gate_120(G352gat,muxed162,G304gat);
nand gate_121(G353gat,G337gat,G305gat);
nand gate_122(G354gat,G339gat,muxed20);
nand gate_123(G355gat,G341gat,muxed149);
nand gate_124(G356gat,muxed135,muxed141);
and gate_125(G357gat,muxed13,muxed8,muxed46,G351gat,muxed161,G353gat,muxed18,muxed148,muxed131);
not gate_126(G360gat,muxed15);
not gate_127(G370gat,muxed15);
nand gate_128(G371gat,G14gat,muxed120);
nand gate_129(G372gat,muxed120,G27gat);
nand gate_130(G373gat,muxed120,G40gat);
nand gate_131(G374gat,muxed120,G53gat);
nand gate_132(G375gat,muxed120,G66gat);
nand gate_133(G376gat,muxed120,G79gat);
nand gate_134(G377gat,muxed120,G92gat);
nand gate_135(G378gat,muxed120,G105gat);
nand gate_136(G379gat,muxed120,G115gat);
nand gate_137(G380gat,G4gat,G242gat,G334gat,G371gat);
nand gate_138(G381gat,muxed99,G336gat,G372gat,G17gat);
nand gate_139(G386gat,muxed93,G338gat,muxed111,G30gat);
nand gate_140(G393gat,G254gat,G340gat,G374gat,muxed189);
nand gate_141(G399gat,muxed65,G342gat,G375gat,G56gat);
nand gate_142(G404gat,muxed184,G344gat,muxed157,G69gat);
nand gate_143(G407gat,G257gat,G345gat,G377gat,G82gat);
nand gate_144(G411gat,G258gat,muxed198,G378gat,G95gat);
nand gate_145(G414gat,G259gat,G347gat,muxed4,G108gat);
not gate_146(G415gat,G380gat);
and gate_147(G416gat,muxed98,muxed176,G393gat,G399gat,muxed152,G407gat,muxed85,muxed2);
not gate_148(G417gat,G393gat);
not gate_149(G418gat,muxed152);
not gate_150(G419gat,G407gat);
not gate_151(G420gat,muxed85);
nor gate_152(G421gat,G415gat,muxed102);
nand gate_153(G422gat,muxed176,G417gat);
nand gate_154(G425gat,muxed176,G393gat,G418gat,G399gat);
nand gate_155(G428gat,G399gat,G393gat,muxed53);
nand gate_156(G429gat,muxed176,G393gat,G407gat,G420gat);
nand gate_157(G430gat,muxed98,muxed176,G422gat,G399gat);
nand gate_158(G431gat,muxed98,muxed176,muxed187,muxed49);
nand gate_159(G432gat,muxed98,G422gat,muxed187,G429gat);
assign muxed0 = keyinput0 ? muxed9 : muxed102;
assign muxed1 = keyinput1 ? muxed96 : muxed83;
assign muxed2 = keyinput2 ? G414gat : muxed32;
assign muxed3 = keyinput3 ? G146gat : G414gat;
assign muxed4 = keyinput4 ? muxed166 : G375gat;
assign muxed5 = keyinput5 ? G184gat : muxed166;
assign muxed6 = keyinput6 ? G360gat : muxed123;
assign muxed7 = keyinput7 ? muxed160 : G185gat;
assign muxed8 = keyinput8 ? G349gat : G377gat;
assign muxed9 = keyinput9 ? G227gat : G349gat;
assign muxed10 = keyinput10 ? muxed60 : muxed141;
assign muxed11 = keyinput11 ? G276gat : muxed60;
assign muxed12 = keyinput12 ? G288gat : G134gat;
assign muxed13 = keyinput13 ? G348gat : G288gat;
assign muxed14 = keyinput14 ? G76gat : muxed15;
assign muxed15 = keyinput15 ? muxed7 : G348gat;
assign muxed16 = keyinput16 ? muxed174 : muxed152;
assign muxed17 = keyinput17 ? muxed52 : muxed174;
assign muxed18 = keyinput18 ? G354gat : muxed166;
assign muxed19 = keyinput19 ? muxed87 : G354gat;
assign muxed20 = keyinput20 ? G306gat : G165gat;
assign muxed21 = keyinput21 ? G331gat : G306gat;
assign muxed22 = keyinput22 ? muxed190 : G341gat;
assign muxed23 = keyinput23 ? G282gat : muxed190;
assign muxed24 = keyinput24 ? muxed31 : G168gat;
assign muxed25 = keyinput25 ? muxed59 : G377gat;
assign muxed26 = keyinput26 ? G142gat : muxed38;
assign muxed27 = keyinput27 ? G119gat : G142gat;
assign muxed28 = keyinput28 ? G43gat : muxed190;
assign muxed29 = keyinput29 ? muxed76 : muxed191;
assign muxed30 = keyinput30 ? muxed24 : G171gat;
assign muxed31 = keyinput31 ? G243gat : G168gat;
assign muxed32 = keyinput32 ? G127gat : G243gat;
assign muxed33 = keyinput33 ? muxed56 : G377gat;
assign muxed34 = keyinput34 ? G174gat : muxed160;
assign muxed35 = keyinput35 ? G236gat : G174gat;
assign muxed36 = keyinput36 ? muxed132 : G142gat;
assign muxed37 = keyinput37 ? muxed133 : muxed132;
assign muxed38 = keyinput38 ? muxed172 : muxed170;
assign muxed39 = keyinput39 ? G131gat : G353gat;
assign muxed40 = keyinput40 ? muxed173 : muxed56;
assign muxed41 = keyinput41 ? muxed57 : G417gat;
assign muxed42 = keyinput42 ? muxed159 : muxed100;
assign muxed43 = keyinput43 ? G376gat : muxed159;
assign muxed44 = keyinput44 ? muxed67 : muxed161;
assign muxed45 = keyinput45 ? muxed145 : G192gat;
assign muxed46 = keyinput46 ? muxed69 : muxed148;
assign muxed47 = keyinput47 ? muxed197 : muxed69;
assign muxed48 = keyinput48 ? G302gat : muxed102;
assign muxed49 = keyinput49 ? muxed58 : G302gat;
assign muxed50 = keyinput50 ? muxed144 : muxed187;
assign muxed51 = keyinput51 ? muxed106 : muxed144;
assign muxed52 = keyinput52 ? G289gat : muxed13;
assign muxed53 = keyinput53 ? muxed107 : G289gat;
assign muxed54 = keyinput54 ? G102gat : muxed170;
assign muxed55 = keyinput55 ? muxed171 : G339gat;
assign muxed56 = keyinput56 ? muxed41 : G407gat;
assign muxed57 = keyinput57 ? muxed25 : G127gat;
assign muxed58 = keyinput58 ? G428gat : muxed25;
assign muxed59 = keyinput59 ? muxed42 : muxed12;
assign muxed60 = keyinput60 ? G301gat : muxed42;
assign muxed61 = keyinput61 ? G295gat : muxed65;
assign muxed62 = keyinput62 ? G251gat : muxed22;
assign muxed63 = keyinput63 ? G180gat : G279gat;
assign muxed64 = keyinput64 ? G150gat : muxed32;
assign muxed65 = keyinput65 ? G255gat : G150gat;
assign muxed66 = keyinput66 ? G8gat : muxed67;
assign muxed67 = keyinput67 ? muxed16 : muxed35;
assign muxed68 = keyinput68 ? muxed153 : muxed76;
assign muxed69 = keyinput69 ? G350gat : muxed164;
assign muxed70 = keyinput70 ? muxed79 : muxed56;
assign muxed71 = keyinput71 ? muxed177 : muxed79;
assign muxed72 = keyinput72 ? muxed81 : G194gat;
assign muxed73 = keyinput73 ? muxed84 : G377gat;
assign muxed74 = keyinput74 ? G260gat : muxed87;
assign muxed75 = keyinput75 ? G157gat : muxed52;
assign muxed76 = keyinput76 ? G293gat : G157gat;
assign muxed77 = keyinput77 ? G233gat : muxed166;
assign muxed78 = keyinput78 ? muxed116 : muxed145;
assign muxed79 = keyinput79 ? muxed48 : muxed174;
assign muxed80 = keyinput80 ? muxed103 : muxed41;
assign muxed81 = keyinput81 ? muxed95 : G422gat;
assign muxed82 = keyinput82 ? G135gat : muxed95;
assign muxed83 = keyinput83 ? muxed73 : G351gat;
assign muxed84 = keyinput84 ? G330gat : G414gat;
assign muxed85 = keyinput85 ? G411gat : G330gat;
assign muxed86 = keyinput86 ? muxed74 : muxed7;
assign muxed87 = keyinput87 ? G290gat : muxed176;
assign muxed88 = keyinput88 ? G213gat : muxed178;
assign muxed89 = keyinput89 ? muxed179 : G376gat;
assign muxed90 = keyinput90 ? muxed105 : G127gat;
assign muxed91 = keyinput91 ? muxed72 : muxed105;
assign muxed92 = keyinput92 ? muxed108 : muxed187;
assign muxed93 = keyinput93 ? muxed136 : muxed108;
assign muxed94 = keyinput94 ? muxed82 : muxed176;
assign muxed95 = keyinput95 ? muxed193 : muxed49;
assign muxed96 = keyinput96 ? G416gat : G185gat;
assign muxed97 = keyinput97 ? muxed163 : G416gat;
assign muxed98 = keyinput98 ? G381gat : G302gat;
assign muxed99 = keyinput99 ? G246gat : G233gat;
assign muxed100 = keyinput100 ? muxed61 : G246gat;
assign muxed101 = keyinput101 ? muxed121 : muxed102;
assign muxed102 = keyinput102 ? muxed80 : G192gat;
assign muxed103 = keyinput103 ? muxed91 : G194gat;
assign muxed104 = keyinput104 ? G158gat : muxed91;
assign muxed105 = keyinput105 ? muxed51 : muxed88;
assign muxed106 = keyinput106 ? muxed92 : muxed178;
assign muxed107 = keyinput107 ? G419gat : muxed92;
assign muxed108 = keyinput108 ? G190gat : G199gat;
assign muxed109 = keyinput109 ? muxed94 : muxed41;
assign muxed110 = keyinput110 ? G386gat : muxed39;
assign muxed111 = keyinput111 ? G373gat : muxed27;
assign muxed112 = keyinput112 ? muxed181 : G373gat;
assign muxed113 = keyinput113 ? muxed86 : muxed114;
assign muxed114 = keyinput114 ? muxed126 : muxed80;
assign muxed115 = keyinput115 ? muxed128 : muxed186;
assign muxed116 = keyinput116 ? muxed139 : G276gat;
assign muxed117 = keyinput117 ? G250gat : muxed139;
assign muxed118 = keyinput118 ? G379gat : muxed7;
assign muxed119 = keyinput119 ? G126gat : G379gat;
assign muxed120 = keyinput120 ? muxed101 : muxed5;
assign muxed121 = keyinput121 ? muxed6 : muxed6;
assign muxed122 = keyinput122 ? muxed64 : muxed6;
assign muxed123 = keyinput123 ? G319gat : muxed193;
assign muxed124 = keyinput124 ? G296gat : muxed73;
assign muxed125 = keyinput125 ? muxed62 : muxed126;
assign muxed126 = keyinput126 ? muxed165 : muxed65;
assign muxed127 = keyinput127 ? muxed167 : muxed108;
assign muxed128 = keyinput128 ? muxed156 : muxed136;
assign muxed129 = keyinput129 ? muxed118 : muxed156;
assign muxed130 = keyinput130 ? muxed146 : muxed49;
assign muxed131 = keyinput131 ? muxed37 : muxed48;
assign muxed132 = keyinput132 ? muxed26 : muxed37;
assign muxed133 = keyinput133 ? G356gat : muxed65;
assign muxed134 = keyinput134 ? muxed143 : G356gat;
assign muxed135 = keyinput135 ? G343gat : G185gat;
assign muxed136 = keyinput136 ? muxed117 : G343gat;
assign muxed137 = keyinput137 ? muxed150 : G341gat;
assign muxed138 = keyinput138 ? G294gat : muxed139;
assign muxed139 = keyinput139 ? muxed71 : muxed109;
assign muxed140 = keyinput140 ? muxed129 : muxed178;
assign muxed141 = keyinput141 ? G308gat : muxed129;
assign muxed142 = keyinput142 ? muxed134 : G260gat;
assign muxed143 = keyinput143 ? muxed78 : G381gat;
assign muxed144 = keyinput144 ? muxed17 : muxed78;
assign muxed145 = keyinput145 ? muxed130 : muxed38;
assign muxed146 = keyinput146 ? G357gat : G146gat;
assign muxed147 = keyinput147 ? G197gat : G357gat;
assign muxed148 = keyinput148 ? G355gat : muxed93;
assign muxed149 = keyinput149 ? G307gat : muxed124;
assign muxed150 = keyinput150 ? G285gat : G307gat;
assign muxed151 = keyinput151 ? G309gat : muxed152;
assign muxed152 = keyinput152 ? muxed68 : muxed145;
assign muxed153 = keyinput153 ? muxed196 : G422gat;
assign muxed154 = keyinput154 ? muxed104 : muxed196;
assign muxed155 = keyinput155 ? G404gat : muxed199;
assign muxed156 = keyinput156 ? muxed142 : G404gat;
assign muxed157 = keyinput157 ? muxed43 : muxed87;
assign muxed158 = keyinput158 ? G122gat : muxed43;
assign muxed159 = keyinput159 ? muxed34 : muxed81;
assign muxed160 = keyinput160 ? muxed44 : G393gat;
assign muxed161 = keyinput161 ? G352gat : muxed67;
assign muxed162 = keyinput162 ? muxed182 : G373gat;
assign muxed163 = keyinput163 ? G159gat : muxed182;
assign muxed164 = keyinput164 ? muxed119 : muxed165;
assign muxed165 = keyinput165 ? muxed77 : G393gat;
assign muxed166 = keyinput166 ? muxed127 : G123gat;
assign muxed167 = keyinput167 ? muxed185 : muxed26;
assign muxed168 = keyinput168 ? muxed90 : muxed185;
assign muxed169 = keyinput169 ? muxed54 : muxed187;
assign muxed170 = keyinput170 ? muxed55 : G122gat;
assign muxed171 = keyinput171 ? muxed40 : muxed72;
assign muxed172 = keyinput172 ? G188gat : muxed40;
assign muxed173 = keyinput173 ? G230gat : muxed85;
assign muxed174 = keyinput174 ? muxed45 : G230gat;
assign muxed175 = keyinput175 ? G162gat : G330gat;
assign muxed176 = keyinput176 ? muxed110 : muxed177;
assign muxed177 = keyinput177 ? muxed140 : G254gat;
assign muxed178 = keyinput178 ? muxed195 : G267gat;
assign muxed179 = keyinput179 ? muxed112 : G307gat;
assign muxed180 = keyinput180 ? G193gat : muxed112;
assign muxed181 = keyinput181 ? G291gat : muxed14;
assign muxed182 = keyinput182 ? G335gat : G291gat;
assign muxed183 = keyinput183 ? muxed168 : muxed161;
assign muxed184 = keyinput184 ? G256gat : muxed168;
assign muxed185 = keyinput185 ? muxed115 : muxed114;
assign muxed186 = keyinput186 ? muxed169 : G242gat;
assign muxed187 = keyinput187 ? G425gat : muxed161;
assign muxed188 = keyinput188 ? G239gat : muxed189;
assign muxed189 = keyinput189 ? muxed28 : G251gat;
assign muxed190 = keyinput190 ? muxed29 : muxed86;
assign muxed191 = keyinput191 ? G300gat : muxed93;
assign muxed192 = keyinput192 ? G263gat : muxed83;
assign muxed193 = keyinput193 ? muxed1 : G263gat;
assign muxed194 = keyinput194 ? muxed154 : G177gat;
assign muxed195 = keyinput195 ? muxed89 : muxed154;
assign muxed196 = keyinput196 ? muxed47 : G332gat;
assign muxed197 = keyinput197 ? muxed155 : G158gat;
assign muxed198 = keyinput198 ? G346gat : muxed155;
assign muxed199 = keyinput199 ? G292gat : G425gat;
endmodule
