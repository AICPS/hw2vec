`timescale 1ns / 1ps
module top (G1,G10,G11,G12,G13,G1324,G1325,G1326,G1327,G1328,G1329,G1330,
  G1331,G1332,G1333,G1334,G1335,G1336,G1337,G1338,G1339,G1340,G1341,G1342,
  G1343,G1344,G1345,G1346,G1347,G1348,G1349,G1350,G1351,G1352,G1353,G1354,
  G1355,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G3,
                  G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G4,G40,G41,G5,G6,G7,G8,G9,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
        keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
                  keyinput125, keyinput126, keyinput127,
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202,
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207,
                  keyinput208, keyinput209,
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
        keyinput250);

  input keyinput210, keyinput211, keyinput212, keyinput213, keyinput214;
  input keyinput215, keyinput216, keyinput217, keyinput218, keyinput219;
  input keyinput220, keyinput221, keyinput222, keyinput223, keyinput224;
  input keyinput225, keyinput226, keyinput227, keyinput228, keyinput229;
  input keyinput230, keyinput231, keyinput232, keyinput233, keyinput234;
  input keyinput235, keyinput236, keyinput237, keyinput238, keyinput239;
  input keyinput240, keyinput241, keyinput242, keyinput243, keyinput244;
  input keyinput245, keyinput246, keyinput247, keyinput248, keyinput249;
  input keyinput250;


  input keyinput128, keyinput129, keyinput130, keyinput131, keyinput132;
  input keyinput133, keyinput134, keyinput135, keyinput136, keyinput137;
  input keyinput138, keyinput139, keyinput140, keyinput141, keyinput142;
  input keyinput143, keyinput144, keyinput145, keyinput146, keyinput147;
  input keyinput148, keyinput149, keyinput150, keyinput151, keyinput152;
  input keyinput153, keyinput154, keyinput155, keyinput156, keyinput157;
  input keyinput158, keyinput159, keyinput160, keyinput161, keyinput162;
  input keyinput163, keyinput164, keyinput165, keyinput166, keyinput167;
  input keyinput168, keyinput169, keyinput170, keyinput171, keyinput172;
  input keyinput173, keyinput174, keyinput175, keyinput176, keyinput177;
  input keyinput178, keyinput179, keyinput180, keyinput181, keyinput182;
  input keyinput183, keyinput184, keyinput185, keyinput186, keyinput187;
  input keyinput188, keyinput189, keyinput190, keyinput191, keyinput192;
  input keyinput193, keyinput194, keyinput195, keyinput196, keyinput197;
  input keyinput198, keyinput199, keyinput200, keyinput201, keyinput202;
  input keyinput203, keyinput204, keyinput205, keyinput206, keyinput207;
  input keyinput208, keyinput209;

  wire KeyWire_0_1 , KeyWire_0_2;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31, keyinput32, keyinput33, keyinput34;
  input keyinput35, keyinput36, keyinput37, keyinput38, keyinput39;
  input keyinput40, keyinput41, keyinput42, keyinput43, keyinput44;
  input keyinput45, keyinput46, keyinput47, keyinput48, keyinput49;
  input keyinput50, keyinput51, keyinput52, keyinput53, keyinput54;
  input keyinput55, keyinput56, keyinput57, keyinput58, keyinput59;
  input keyinput60, keyinput61, keyinput62, keyinput63, keyinput64;
  input keyinput65, keyinput66, keyinput67, keyinput68, keyinput69;
  input keyinput70, keyinput71, keyinput72, keyinput73, keyinput74;
  input keyinput75, keyinput76, keyinput77, keyinput78, keyinput79;
  input keyinput80, keyinput81, keyinput82, keyinput83, keyinput84;
  input keyinput85, keyinput86, keyinput87, keyinput88, keyinput89;
  input keyinput90, keyinput91, keyinput92, keyinput93, keyinput94;
  input keyinput95, keyinput96, keyinput97, keyinput98, keyinput99;
  input keyinput100, keyinput101, keyinput102, keyinput103, keyinput104;
  input keyinput105, keyinput106, keyinput107, keyinput108, keyinput109;
  input keyinput110, keyinput111, keyinput112, keyinput113, keyinput114;
  input keyinput115, keyinput116, keyinput117, keyinput118, keyinput119;
  input keyinput120, keyinput121, keyinput122, keyinput123, keyinput124;
  input keyinput125, keyinput126, keyinput127;

  wire [0:127] keyinput_Wire_0;
  wire [0:64] KeyNOTWire_0;
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
  G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,
  G40,G41;
output G1324,G1325,G1326,G1327,G1328,G1329,G1330,G1331,G1332,G1333,G1334,G1335,
  G1336,G1337,G1338,G1339,G1340,G1341,G1342,G1343,G1344,G1345,G1346,G1347,
  G1348,G1349,G1350,G1351,G1352,G1353,G1354,G1355;

  wire G242,G245,G248,G251,G254,G257,G260,G263,G266,G269,G272,G275,G278,G281,
    G284,G287,G290,G293,G296,G299,G302,G305,G308,G311,G314,G317,G320,G323,G326,
    G329,G332,G335,G338,G341,G344,G347,G350,G353,G356,G359,G362,G363,G364,G365,
    G366,G367,G368,G369,G370,G371,G372,G373,G374,G375,G376,G377,G378,G379,G380,
    G381,G382,G383,G384,G385,G386,G387,G388,G389,G390,G391,G392,G393,G394,G395,
    G396,G397,G398,G399,G400,G401,G402,G403,G404,G405,G406,G407,G408,G409,G410,
    G411,G412,G413,G414,G415,G416,G417,G418,G419,G420,G421,G422,G423,G424,G425,
    G426,G429,G432,G435,G438,G441,G444,G447,G450,G453,G456,G459,G462,G465,G468,
    G471,G474,G477,G480,G483,G486,G489,G492,G495,G498,G501,G504,G507,G510,G513,
    G516,G519,G522,G525,G528,G531,G534,G537,G540,G543,G546,G549,G552,G555,G558,
    G561,G564,G567,G570,G571,G572,G573,G574,G575,G576,G577,G578,G579,G580,G581,
    G582,G583,G584,G585,G586,G587,G588,G589,G590,G591,G592,G593,G594,G595,G596,
    G597,G598,G599,G600,G601,G602,G607,G612,G617,G622,G627,G632,G637,G642,G645,
    G648,G651,G654,G657,G660,G663,G666,G669,G672,G675,G678,G681,G684,G687,G690,
    G691,G692,G693,G694,G695,G696,G697,G698,G699,G700,G701,G702,G703,G704,G705,
    G706,G709,G712,G715,G718,G721,G724,G727,G730,G733,G736,G739,G742,G745,G748,
    G751,G754,G755,G756,G757,G758,G759,G760,G761,G762,G763,G764,G765,G766,G767,
    G768,G769,G770,G773,G776,G779,G782,G785,G788,G791,G794,G797,G800,G803,G806,
    G809,G812,G815,G818,G819,G820,G821,G822,G823,G824,G825,G826,G827,G828,G829,
    G830,G831,G832,G833,G834,G847,G860,G873,G886,G899,G912,G925,G938,G939,G940,
    G941,G942,G943,G944,G945,G946,G947,G948,G949,G950,G951,G952,G953,G954,G955,
    G956,G957,G958,G959,G960,G961,G962,G963,G964,G965,G966,G967,G968,G969,G970,
    G971,G972,G973,G974,G975,G976,G977,G978,G979,G980,G981,G982,G983,G984,G985,
    G986,G991,G996,G1001,G1006,G1011,G1016,G1021,G1026,G1031,G1036,G1039,G1042,
    G1045,G1048,G1051,G1054,G1057,G1060,G1063,G1066,G1069,G1072,G1075,G1078,
    G1081,G1084,G1087,G1090,G1093,G1096,G1099,G1102,G1105,G1108,G1111,G1114,
    G1117,G1120,G1123,G1126,G1129,G1132,G1135,G1138,G1141,G1144,G1147,G1150,
    G1153,G1156,G1159,G1162,G1165,G1168,G1171,G1174,G1177,G1180,G1183,G1186,
    G1189,G1192,G1195,G1198,G1201,G1204,G1207,G1210,G1213,G1216,G1219,G1222,
    G1225,G1228,G1229,G1230,G1231,G1232,G1233,G1234,G1235,G1236,G1237,G1238,
    G1239,G1240,G1241,G1242,G1243,G1244,G1245,G1246,G1247,G1248,G1249,G1250,
    G1251,G1252,G1253,G1254,G1255,G1256,G1257,G1258,G1259,G1260,G1261,G1262,
    G1263,G1264,G1265,G1266,G1267,G1268,G1269,G1270,G1271,G1272,G1273,G1274,
    G1275,G1276,G1277,G1278,G1279,G1280,G1281,G1282,G1283,G1284,G1285,G1286,
    G1287,G1288,G1289,G1290,G1291,G1292,G1293,G1294,G1295,G1296,G1297,G1298,
    G1299,G1300,G1301,G1302,G1303,G1304,G1305,G1306,G1307,G1308,G1309,G1310,
    G1311,G1312,G1313,G1314,G1315,G1316,G1317,G1318,G1319,G1320,G1321,G1322,
    G1323;

  and AND2_0(keyinput_Wire_0[0], G33,G41);
  xnor keyGate_0_0(G242, keyinput0, keyinput_Wire_0[0]);
  and AND2_1(keyinput_Wire_0[1], G34,G41);
  xnor keyGate_0_1(G245, keyinput1, keyinput_Wire_0[1]);
  and AND2_2(keyinput_Wire_0[2], G35,G41);
  xor keyGate_0_2(G248, keyinput2, keyinput_Wire_0[2]);
  and AND2_3(G251,G36,G41);
  and AND2_4(keyinput_Wire_0[3], G37,G41);
  xnor keyGate_0_3(KeyNOTWire_0[0], keyinput3, keyinput_Wire_0[3]);
  not KeyNOTGate_0_0(G254, KeyNOTWire_0[0]);
  and AND2_5(G257,G38,G41);
  and AND2_6(keyinput_Wire_0[4], G39,G41);
  xnor keyGate_0_4(KeyNOTWire_0[1], keyinput4, keyinput_Wire_0[4]);
  not KeyNOTGate_0_1(G260, KeyNOTWire_0[1]);
  and AND2_7(G263,G40,G41);
  nand NAND2_0(keyinput_Wire_0[5], G1,G2);
  xor keyGate_0_5(G266, keyinput5, keyinput_Wire_0[5]);
  nand NAND2_1(G269,G3,G4);
  nand NAND2_2(G272,G5,G6);
  nand NAND2_3(G275,G7,G8);
  nand NAND2_4(G278,G9,G10);
  nand NAND2_5(G281,G11,G12);
  nand NAND2_6(keyinput_Wire_0[6], G13,G14);
  xnor keyGate_0_6(G284, keyinput6, keyinput_Wire_0[6]);
  nand NAND2_7(G287,G15,G16);
  nand NAND2_8(keyinput_Wire_0[7], G17,G18);
  xnor keyGate_0_7(G290, keyinput7, keyinput_Wire_0[7]);
  nand NAND2_9(keyinput_Wire_0[8], G19,G20);
  xnor keyGate_0_8(G293, keyinput8, keyinput_Wire_0[8]);
  nand NAND2_10(G296,G21,G22);
  nand NAND2_11(G299,G23,G24);
  nand NAND2_12(G302,G25,G26);
  nand NAND2_13(keyinput_Wire_0[9], G27,G28);
  xnor keyGate_0_9(G305, keyinput9, keyinput_Wire_0[9]);
  nand NAND2_14(G308,G29,G30);
  nand NAND2_15(keyinput_Wire_0[10], G31,G32);
  xor keyGate_0_10(KeyNOTWire_0[2], keyinput10, keyinput_Wire_0[10]);
  not KeyNOTGate_0_2(G311, KeyNOTWire_0[2]);
  nand NAND2_16(G314,G1,G5);
  nand NAND2_17(keyinput_Wire_0[11], G9,G13);
  xor keyGate_0_11(G317, keyinput11, keyinput_Wire_0[11]);
  nand NAND2_18(G320,G2,G6);
  nand NAND2_19(G323,G10,G14);
  nand NAND2_20(G326,G3,G7);
  nand NAND2_21(G329,G11,G15);
  nand NAND2_22(G332,G4,G8);
  nand NAND2_23(G335,G12,G16);
  nand NAND2_24(G338,G17,G21);
  nand NAND2_25(G341,G25,G29);
  nand NAND2_26(keyinput_Wire_0[12], G18,G22);
  xnor keyGate_0_12(G344, keyinput12, keyinput_Wire_0[12]);
  nand NAND2_27(keyinput_Wire_0[13], G26,G30);
  xnor keyGate_0_13(G347, keyinput13, keyinput_Wire_0[13]);
  nand NAND2_28(keyinput_Wire_0[14], G19,G23);
  xor keyGate_0_14(KeyNOTWire_0[3], keyinput14, keyinput_Wire_0[14]);
  not KeyNOTGate_0_3(G350, KeyNOTWire_0[3]);
  nand NAND2_29(G353,G27,G31);
  nand NAND2_30(G356,G20,G24);
  nand NAND2_31(G359,G28,G32);
  nand NAND2_32(keyinput_Wire_0[15], G1,G266);
  xnor keyGate_0_15(G362, keyinput15, keyinput_Wire_0[15]);
  nand NAND2_33(keyinput_Wire_0[16], G2,G266);
  xnor keyGate_0_16(G363, keyinput16, keyinput_Wire_0[16]);
  nand NAND2_34(G364,G3,G269);
  nand NAND2_35(G365,G4,G269);
  nand NAND2_36(keyinput_Wire_0[17], G5,G272);
  xnor keyGate_0_17(G366, keyinput17, keyinput_Wire_0[17]);
  nand NAND2_37(G367,G6,G272);
  nand NAND2_38(keyinput_Wire_0[18], G7,G275);
  xor keyGate_0_18(G368, keyinput18, keyinput_Wire_0[18]);
  nand NAND2_39(G369,G8,G275);
  nand NAND2_40(G370,G9,G278);
  nand NAND2_41(keyinput_Wire_0[19], G10,G278);
  xnor keyGate_0_19(G371, keyinput19, keyinput_Wire_0[19]);
  nand NAND2_42(G372,G11,G281);
  nand NAND2_43(G373,G12,G281);
  nand NAND2_44(keyinput_Wire_0[20], G13,G284);
  xor keyGate_0_20(G374, keyinput20, keyinput_Wire_0[20]);
  nand NAND2_45(keyinput_Wire_0[21], G14,G284);
  xnor keyGate_0_21(G375, keyinput21, keyinput_Wire_0[21]);
  nand NAND2_46(keyinput_Wire_0[22], G15,G287);
  xor keyGate_0_22(KeyNOTWire_0[4], keyinput22, keyinput_Wire_0[22]);
  not KeyNOTGate_0_4(G376, KeyNOTWire_0[4]);
  nand NAND2_47(keyinput_Wire_0[23], G16,G287);
  xnor keyGate_0_23(KeyNOTWire_0[5], keyinput23, keyinput_Wire_0[23]);
  not KeyNOTGate_0_5(G377, KeyNOTWire_0[5]);
  nand NAND2_48(G378,G17,G290);
  nand NAND2_49(keyinput_Wire_0[24], G18,G290);
  xor keyGate_0_24(G379, keyinput24, keyinput_Wire_0[24]);
  nand NAND2_50(G380,G19,G293);
  nand NAND2_51(keyinput_Wire_0[25], G20,G293);
  xor keyGate_0_25(G381, keyinput25, keyinput_Wire_0[25]);
  nand NAND2_52(G382,G21,G296);
  nand NAND2_53(keyinput_Wire_0[26], G22,G296);
  xnor keyGate_0_26(KeyNOTWire_0[6], keyinput26, keyinput_Wire_0[26]);
  not KeyNOTGate_0_6(G383, KeyNOTWire_0[6]);
  nand NAND2_54(G384,G23,G299);
  nand NAND2_55(G385,G24,G299);
  nand NAND2_56(G386,G25,G302);
  nand NAND2_57(keyinput_Wire_0[27], G26,G302);
  xor keyGate_0_27(KeyNOTWire_0[7], keyinput27, keyinput_Wire_0[27]);
  not KeyNOTGate_0_7(G387, KeyNOTWire_0[7]);
  nand NAND2_58(G388,G27,G305);
  nand NAND2_59(keyinput_Wire_0[28], G28,G305);
  xor keyGate_0_28(G389, keyinput28, keyinput_Wire_0[28]);
  nand NAND2_60(G390,G29,G308);
  nand NAND2_61(keyinput_Wire_0[29], G30,G308);
  xor keyGate_0_29(KeyNOTWire_0[8], keyinput29, keyinput_Wire_0[29]);
  not KeyNOTGate_0_8(G391, KeyNOTWire_0[8]);
  nand NAND2_62(G392,G31,G311);
  nand NAND2_63(keyinput_Wire_0[30], G32,G311);
  xor keyGate_0_30(KeyNOTWire_0[9], keyinput30, keyinput_Wire_0[30]);
  not KeyNOTGate_0_9(G393, KeyNOTWire_0[9]);
  nand NAND2_64(G394,G1,G314);
  nand NAND2_65(G395,G5,G314);
  nand NAND2_66(G396,G9,G317);
  nand NAND2_67(keyinput_Wire_0[31], G13,G317);
  xor keyGate_0_31(KeyNOTWire_0[10], keyinput31, keyinput_Wire_0[31]);
  not KeyNOTGate_0_10(G397, KeyNOTWire_0[10]);
  nand NAND2_68(G398,G2,G320);
  nand NAND2_69(G399,G6,G320);
  nand NAND2_70(G400,G10,G323);
  nand NAND2_71(G401,G14,G323);
  nand NAND2_72(G402,G3,G326);
  nand NAND2_73(G403,G7,G326);
  nand NAND2_74(keyinput_Wire_0[32], G11,G329);
  xnor keyGate_0_32(G404, keyinput32, keyinput_Wire_0[32]);
  nand NAND2_75(G405,G15,G329);
  nand NAND2_76(G406,G4,G332);
  nand NAND2_77(G407,G8,G332);
  nand NAND2_78(G408,G12,G335);
  nand NAND2_79(keyinput_Wire_0[33], G16,G335);
  xnor keyGate_0_33(KeyNOTWire_0[11], keyinput33, keyinput_Wire_0[33]);
  not KeyNOTGate_0_11(G409, KeyNOTWire_0[11]);
  nand NAND2_80(G410,G17,G338);
  nand NAND2_81(G411,G21,G338);
  nand NAND2_82(keyinput_Wire_0[34], G25,G341);
  xnor keyGate_0_34(G412, keyinput34, keyinput_Wire_0[34]);
  nand NAND2_83(G413,G29,G341);
  nand NAND2_84(G414,G18,G344);
  nand NAND2_85(keyinput_Wire_0[35], G22,G344);
  xnor keyGate_0_35(G415, keyinput35, keyinput_Wire_0[35]);
  nand NAND2_86(keyinput_Wire_0[36], G26,G347);
  xnor keyGate_0_36(KeyNOTWire_0[12], keyinput36, keyinput_Wire_0[36]);
  not KeyNOTGate_0_12(G416, KeyNOTWire_0[12]);
  nand NAND2_87(keyinput_Wire_0[37], G30,G347);
  xnor keyGate_0_37(KeyNOTWire_0[13], keyinput37, keyinput_Wire_0[37]);
  not KeyNOTGate_0_13(G417, KeyNOTWire_0[13]);
  nand NAND2_88(G418,G19,G350);
  nand NAND2_89(keyinput_Wire_0[38], G23,G350);
  xor keyGate_0_38(KeyNOTWire_0[14], keyinput38, keyinput_Wire_0[38]);
  not KeyNOTGate_0_14(G419, KeyNOTWire_0[14]);
  nand NAND2_90(G420,G27,G353);
  nand NAND2_91(G421,G31,G353);
  nand NAND2_92(keyinput_Wire_0[39], G20,G356);
  xnor keyGate_0_39(KeyNOTWire_0[15], keyinput39, keyinput_Wire_0[39]);
  not KeyNOTGate_0_15(G422, KeyNOTWire_0[15]);
  nand NAND2_93(G423,G24,G356);
  nand NAND2_94(keyinput_Wire_0[40], G28,G359);
  xor keyGate_0_40(G424, keyinput40, keyinput_Wire_0[40]);
  nand NAND2_95(G425,G32,G359);
  nand NAND2_96(G426,G362,G363);
  nand NAND2_97(G429,G364,G365);
  nand NAND2_98(keyinput_Wire_0[41], G366,G367);
  xor keyGate_0_41(G432, keyinput41, keyinput_Wire_0[41]);
  nand NAND2_99(keyinput_Wire_0[42], G368,G369);
  xor keyGate_0_42(KeyNOTWire_0[16], keyinput42, keyinput_Wire_0[42]);
  not KeyNOTGate_0_16(G435, KeyNOTWire_0[16]);
  nand NAND2_100(keyinput_Wire_0[43], G370,G371);
  xor keyGate_0_43(KeyNOTWire_0[17], keyinput43, keyinput_Wire_0[43]);
  not KeyNOTGate_0_17(G438, KeyNOTWire_0[17]);
  nand NAND2_101(G441,G372,G373);
  nand NAND2_102(G444,G374,G375);
  nand NAND2_103(keyinput_Wire_0[44], G376,G377);
  xor keyGate_0_44(KeyNOTWire_0[18], keyinput44, keyinput_Wire_0[44]);
  not KeyNOTGate_0_18(G447, KeyNOTWire_0[18]);
  nand NAND2_104(G450,G378,G379);
  nand NAND2_105(keyinput_Wire_0[45], G380,G381);
  xnor keyGate_0_45(G453, keyinput45, keyinput_Wire_0[45]);
  nand NAND2_106(G456,G382,G383);
  nand NAND2_107(G459,G384,G385);
  nand NAND2_108(G462,G386,G387);
  nand NAND2_109(G465,G388,G389);
  nand NAND2_110(keyinput_Wire_0[46], G390,G391);
  xnor keyGate_0_46(KeyNOTWire_0[19], keyinput46, keyinput_Wire_0[46]);
  not KeyNOTGate_0_19(G468, KeyNOTWire_0[19]);
  nand NAND2_111(G471,G392,G393);
  nand NAND2_112(keyinput_Wire_0[47], G394,G395);
  xnor keyGate_0_47(G474, keyinput47, keyinput_Wire_0[47]);
  nand NAND2_113(G477,G396,G397);
  nand NAND2_114(keyinput_Wire_0[48], G398,G399);
  xor keyGate_0_48(KeyNOTWire_0[20], keyinput48, keyinput_Wire_0[48]);
  not KeyNOTGate_0_20(G480, KeyNOTWire_0[20]);
  nand NAND2_115(keyinput_Wire_0[49], G400,G401);
  xnor keyGate_0_49(KeyNOTWire_0[21], keyinput49, keyinput_Wire_0[49]);
  not KeyNOTGate_0_21(G483, KeyNOTWire_0[21]);
  nand NAND2_116(keyinput_Wire_0[50], G402,G403);
  xnor keyGate_0_50(KeyNOTWire_0[22], keyinput50, keyinput_Wire_0[50]);
  not KeyNOTGate_0_22(G486, KeyNOTWire_0[22]);
  nand NAND2_117(G489,G404,G405);
  nand NAND2_118(keyinput_Wire_0[51], G406,G407);
  xor keyGate_0_51(KeyNOTWire_0[23], keyinput51, keyinput_Wire_0[51]);
  not KeyNOTGate_0_23(G492, KeyNOTWire_0[23]);
  nand NAND2_119(G495,G408,G409);
  nand NAND2_120(keyinput_Wire_0[52], G410,G411);
  xor keyGate_0_52(G498, keyinput52, keyinput_Wire_0[52]);
  nand NAND2_121(G501,G412,G413);
  nand NAND2_122(G504,G414,G415);
  nand NAND2_123(G507,G416,G417);
  nand NAND2_124(G510,G418,G419);
  nand NAND2_125(G513,G420,G421);
  nand NAND2_126(G516,G422,G423);
  nand NAND2_127(G519,G424,G425);
  nand NAND2_128(keyinput_Wire_0[53], G426,G429);
  xor keyGate_0_53(KeyNOTWire_0[24], keyinput53, keyinput_Wire_0[53]);
  not KeyNOTGate_0_24(G522, KeyNOTWire_0[24]);
  nand NAND2_129(G525,G432,G435);
  nand NAND2_130(G528,G438,G441);
  nand NAND2_131(G531,G444,G447);
  nand NAND2_132(G534,G450,G453);
  nand NAND2_133(G537,G456,G459);
  nand NAND2_134(keyinput_Wire_0[54], G462,G465);
  xnor keyGate_0_54(G540, keyinput54, keyinput_Wire_0[54]);
  nand NAND2_135(G543,G468,G471);
  nand NAND2_136(G546,G474,G477);
  nand NAND2_137(keyinput_Wire_0[55], G480,G483);
  xor keyGate_0_55(KeyNOTWire_0[25], keyinput55, keyinput_Wire_0[55]);
  not KeyNOTGate_0_25(G549, KeyNOTWire_0[25]);
  nand NAND2_138(G552,G486,G489);
  nand NAND2_139(G555,G492,G495);
  nand NAND2_140(keyinput_Wire_0[56], G498,G501);
  xnor keyGate_0_56(KeyNOTWire_0[26], keyinput56, keyinput_Wire_0[56]);
  not KeyNOTGate_0_26(G558, KeyNOTWire_0[26]);
  nand NAND2_141(keyinput_Wire_0[57], G504,G507);
  xnor keyGate_0_57(KeyNOTWire_0[27], keyinput57, keyinput_Wire_0[57]);
  not KeyNOTGate_0_27(G561, KeyNOTWire_0[27]);
  nand NAND2_142(G564,G510,G513);
  nand NAND2_143(keyinput_Wire_0[58], G516,G519);
  xnor keyGate_0_58(KeyNOTWire_0[28], keyinput58, keyinput_Wire_0[58]);
  not KeyNOTGate_0_28(G567, KeyNOTWire_0[28]);
  nand NAND2_144(G570,G426,G522);
  nand NAND2_145(keyinput_Wire_0[59], G429,G522);
  xor keyGate_0_59(KeyNOTWire_0[29], keyinput59, keyinput_Wire_0[59]);
  not KeyNOTGate_0_29(G571, KeyNOTWire_0[29]);
  nand NAND2_146(keyinput_Wire_0[60], G432,G525);
  xnor keyGate_0_60(G572, keyinput60, keyinput_Wire_0[60]);
  nand NAND2_147(keyinput_Wire_0[61], G435,G525);
  xor keyGate_0_61(KeyNOTWire_0[30], keyinput61, keyinput_Wire_0[61]);
  not KeyNOTGate_0_30(G573, KeyNOTWire_0[30]);
  nand NAND2_148(G574,G438,G528);
  nand NAND2_149(keyinput_Wire_0[62], G441,G528);
  xor keyGate_0_62(G575, keyinput62, keyinput_Wire_0[62]);
  nand NAND2_150(G576,G444,G531);
  nand NAND2_151(G577,G447,G531);
  nand NAND2_152(G578,G450,G534);
  nand NAND2_153(keyinput_Wire_0[63], G453,G534);
  xnor keyGate_0_63(KeyNOTWire_0[31], keyinput63, keyinput_Wire_0[63]);
  not KeyNOTGate_0_31(G579, KeyNOTWire_0[31]);
  nand NAND2_154(keyinput_Wire_0[64], G456,G537);
  xor keyGate_0_64(G580, keyinput64, keyinput_Wire_0[64]);
  nand NAND2_155(G581,G459,G537);
  nand NAND2_156(G582,G462,G540);
  nand NAND2_157(keyinput_Wire_0[65], G465,G540);
  xor keyGate_0_65(G583, keyinput65, keyinput_Wire_0[65]);
  nand NAND2_158(G584,G468,G543);
  nand NAND2_159(G585,G471,G543);
  nand NAND2_160(G586,G474,G546);
  nand NAND2_161(G587,G477,G546);
  nand NAND2_162(G588,G480,G549);
  nand NAND2_163(G589,G483,G549);
  nand NAND2_164(G590,G486,G552);
  nand NAND2_165(keyinput_Wire_0[66], G489,G552);
  xor keyGate_0_66(KeyNOTWire_0[32], keyinput66, keyinput_Wire_0[66]);
  not KeyNOTGate_0_32(G591, KeyNOTWire_0[32]);
  nand NAND2_166(keyinput_Wire_0[67], G492,G555);
  xor keyGate_0_67(KeyNOTWire_0[33], keyinput67, keyinput_Wire_0[67]);
  not KeyNOTGate_0_33(G592, KeyNOTWire_0[33]);
  nand NAND2_167(G593,G495,G555);
  nand NAND2_168(keyinput_Wire_0[68], G498,G558);
  xor keyGate_0_68(G594, keyinput68, keyinput_Wire_0[68]);
  nand NAND2_169(keyinput_Wire_0[69], G501,G558);
  xnor keyGate_0_69(G595, keyinput69, keyinput_Wire_0[69]);
  nand NAND2_170(G596,G504,G561);
  nand NAND2_171(keyinput_Wire_0[70], G507,G561);
  xnor keyGate_0_70(KeyNOTWire_0[34], keyinput70, keyinput_Wire_0[70]);
  not KeyNOTGate_0_34(G597, KeyNOTWire_0[34]);
  nand NAND2_172(G598,G510,G564);
  nand NAND2_173(keyinput_Wire_0[71], G513,G564);
  xor keyGate_0_71(G599, keyinput71, keyinput_Wire_0[71]);
  nand NAND2_174(G600,G516,G567);
  nand NAND2_175(keyinput_Wire_0[72], G519,G567);
  xnor keyGate_0_72(G601, keyinput72, keyinput_Wire_0[72]);
  nand NAND2_176(G602,G570,G571);
  nand NAND2_177(keyinput_Wire_0[73], G572,G573);
  xnor keyGate_0_73(G607, keyinput73, keyinput_Wire_0[73]);
  nand NAND2_178(keyinput_Wire_0[74], G574,G575);
  xor keyGate_0_74(G612, keyinput74, keyinput_Wire_0[74]);
  nand NAND2_179(G617,G576,G577);
  nand NAND2_180(G622,G578,G579);
  nand NAND2_181(G627,G580,G581);
  nand NAND2_182(G632,G582,G583);
  nand NAND2_183(G637,G584,G585);
  nand NAND2_184(keyinput_Wire_0[75], G586,G587);
  xnor keyGate_0_75(KeyNOTWire_0[35], keyinput75, keyinput_Wire_0[75]);
  not KeyNOTGate_0_35(G642, KeyNOTWire_0[35]);
  nand NAND2_185(G645,G588,G589);
  nand NAND2_186(G648,G590,G591);
  nand NAND2_187(G651,G592,G593);
  nand NAND2_188(G654,G594,G595);
  nand NAND2_189(keyinput_Wire_0[76], G596,G597);
  xor keyGate_0_76(KeyNOTWire_0[36], keyinput76, keyinput_Wire_0[76]);
  not KeyNOTGate_0_36(G657, KeyNOTWire_0[36]);
  nand NAND2_190(G660,G598,G599);
  nand NAND2_191(keyinput_Wire_0[77], G600,G601);
  xor keyGate_0_77(G663, keyinput77, keyinput_Wire_0[77]);
  nand NAND2_192(G666,G602,G607);
  nand NAND2_193(G669,G612,G617);
  nand NAND2_194(G672,G602,G612);
  nand NAND2_195(keyinput_Wire_0[78], G607,G617);
  xor keyGate_0_78(G675, keyinput78, keyinput_Wire_0[78]);
  nand NAND2_196(keyinput_Wire_0[79], G622,G627);
  xnor keyGate_0_79(G678, keyinput79, keyinput_Wire_0[79]);
  nand NAND2_197(G681,G632,G637);
  nand NAND2_198(G684,G622,G632);
  nand NAND2_199(keyinput_Wire_0[80], G627,G637);
  xor keyGate_0_80(KeyNOTWire_0[37], keyinput80, keyinput_Wire_0[80]);
  not KeyNOTGate_0_37(G687, KeyNOTWire_0[37]);
  nand NAND2_200(G690,G602,G666);
  nand NAND2_201(keyinput_Wire_0[81], G607,G666);
  xnor keyGate_0_81(G691, keyinput81, keyinput_Wire_0[81]);
  nand NAND2_202(G692,G612,G669);
  nand NAND2_203(G693,G617,G669);
  nand NAND2_204(G694,G602,G672);
  nand NAND2_205(G695,G612,G672);
  nand NAND2_206(G696,G607,G675);
  nand NAND2_207(keyinput_Wire_0[82], G617,G675);
  xor keyGate_0_82(G697, keyinput82, keyinput_Wire_0[82]);
  nand NAND2_208(keyinput_Wire_0[83], G622,G678);
  xnor keyGate_0_83(G698, keyinput83, keyinput_Wire_0[83]);
  nand NAND2_209(keyinput_Wire_0[84], G627,G678);
  xnor keyGate_0_84(KeyNOTWire_0[38], keyinput84, keyinput_Wire_0[84]);
  not KeyNOTGate_0_38(G699, KeyNOTWire_0[38]);
  nand NAND2_210(G700,G632,G681);
  nand NAND2_211(G701,G637,G681);
  nand NAND2_212(G702,G622,G684);
  nand NAND2_213(keyinput_Wire_0[85], G632,G684);
  xnor keyGate_0_85(G703, keyinput85, keyinput_Wire_0[85]);
  nand NAND2_214(G704,G627,G687);
  nand NAND2_215(keyinput_Wire_0[86], G637,G687);
  xnor keyGate_0_86(KeyNOTWire_0[39], keyinput86, keyinput_Wire_0[86]);
  not KeyNOTGate_0_39(G705, KeyNOTWire_0[39]);
  nand NAND2_216(keyinput_Wire_0[87], G690,G691);
  xor keyGate_0_87(KeyNOTWire_0[40], keyinput87, keyinput_Wire_0[87]);
  not KeyNOTGate_0_40(G706, KeyNOTWire_0[40]);
  nand NAND2_217(keyinput_Wire_0[88], G692,G693);
  xor keyGate_0_88(G709, keyinput88, keyinput_Wire_0[88]);
  nand NAND2_218(G712,G694,G695);
  nand NAND2_219(G715,G696,G697);
  nand NAND2_220(G718,G698,G699);
  nand NAND2_221(keyinput_Wire_0[89], G700,G701);
  xor keyGate_0_89(KeyNOTWire_0[41], keyinput89, keyinput_Wire_0[89]);
  not KeyNOTGate_0_41(G721, KeyNOTWire_0[41]);
  nand NAND2_222(G724,G702,G703);
  nand NAND2_223(G727,G704,G705);
  nand NAND2_224(G730,G242,G718);
  nand NAND2_225(keyinput_Wire_0[90], G245,G721);
  xnor keyGate_0_90(KeyNOTWire_0[42], keyinput90, keyinput_Wire_0[90]);
  not KeyNOTGate_0_42(G733, KeyNOTWire_0[42]);
  nand NAND2_226(keyinput_Wire_0[91], G248,G724);
  xor keyGate_0_91(KeyNOTWire_0[43], keyinput91, keyinput_Wire_0[91]);
  not KeyNOTGate_0_43(G736, KeyNOTWire_0[43]);
  nand NAND2_227(keyinput_Wire_0[92], G251,G727);
  xnor keyGate_0_92(KeyNOTWire_0[44], keyinput92, keyinput_Wire_0[92]);
  not KeyNOTGate_0_44(G739, KeyNOTWire_0[44]);
  nand NAND2_228(G742,G254,G706);
  nand NAND2_229(keyinput_Wire_0[93], G257,G709);
  xor keyGate_0_93(KeyNOTWire_0[45], keyinput93, keyinput_Wire_0[93]);
  not KeyNOTGate_0_45(G745, KeyNOTWire_0[45]);
  nand NAND2_230(G748,G260,G712);
  nand NAND2_231(G751,G263,G715);
  nand NAND2_232(G754,G242,G730);
  nand NAND2_233(keyinput_Wire_0[94], G718,G730);
  xor keyGate_0_94(KeyNOTWire_0[46], keyinput94, keyinput_Wire_0[94]);
  not KeyNOTGate_0_46(G755, KeyNOTWire_0[46]);
  nand NAND2_234(G756,G245,G733);
  nand NAND2_235(keyinput_Wire_0[95], G721,G733);
  xnor keyGate_0_95(KeyNOTWire_0[47], keyinput95, keyinput_Wire_0[95]);
  not KeyNOTGate_0_47(G757, KeyNOTWire_0[47]);
  nand NAND2_236(keyinput_Wire_0[96], G248,G736);
  xor keyGate_0_96(G758, keyinput96, keyinput_Wire_0[96]);
  nand NAND2_237(keyinput_Wire_0[97], G724,G736);
  xor keyGate_0_97(KeyNOTWire_0[48], keyinput97, keyinput_Wire_0[97]);
  not KeyNOTGate_0_48(G759, KeyNOTWire_0[48]);
  nand NAND2_238(G760,G251,G739);
  nand NAND2_239(keyinput_Wire_0[98], G727,G739);
  xnor keyGate_0_98(KeyNOTWire_0[49], keyinput98, keyinput_Wire_0[98]);
  not KeyNOTGate_0_49(G761, KeyNOTWire_0[49]);
  nand NAND2_240(G762,G254,G742);
  nand NAND2_241(keyinput_Wire_0[99], G706,G742);
  xor keyGate_0_99(KeyNOTWire_0[50], keyinput99, keyinput_Wire_0[99]);
  not KeyNOTGate_0_50(G763, KeyNOTWire_0[50]);
  nand NAND2_242(keyinput_Wire_0[100], G257,G745);
  xnor keyGate_0_100(KeyNOTWire_0[51], keyinput100, keyinput_Wire_0[100]);
  not KeyNOTGate_0_51(G764, KeyNOTWire_0[51]);
  nand NAND2_243(keyinput_Wire_0[101], G709,G745);
  xor keyGate_0_101(KeyNOTWire_0[52], keyinput101, keyinput_Wire_0[101]);
  not KeyNOTGate_0_52(G765, KeyNOTWire_0[52]);
  nand NAND2_244(G766,G260,G748);
  nand NAND2_245(keyinput_Wire_0[102], G712,G748);
  xor keyGate_0_102(KeyNOTWire_0[53], keyinput102, keyinput_Wire_0[102]);
  not KeyNOTGate_0_53(G767, KeyNOTWire_0[53]);
  nand NAND2_246(G768,G263,G751);
  nand NAND2_247(G769,G715,G751);
  nand NAND2_248(keyinput_Wire_0[103], G754,G755);
  xor keyGate_0_103(G770, keyinput103, keyinput_Wire_0[103]);
  nand NAND2_249(G773,G756,G757);
  nand NAND2_250(keyinput_Wire_0[104], G758,G759);
  xnor keyGate_0_104(G776, keyinput104, keyinput_Wire_0[104]);
  nand NAND2_251(G779,G760,G761);
  nand NAND2_252(keyinput_Wire_0[105], G762,G763);
  xnor keyGate_0_105(KeyNOTWire_0[54], keyinput105, keyinput_Wire_0[105]);
  not KeyNOTGate_0_54(G782, KeyNOTWire_0[54]);
  nand NAND2_253(keyinput_Wire_0[106], G764,G765);
  xnor keyGate_0_106(G785, keyinput106, keyinput_Wire_0[106]);
  nand NAND2_254(G788,G766,G767);
  nand NAND2_255(keyinput_Wire_0[107], G768,G769);
  xor keyGate_0_107(G791, keyinput107, keyinput_Wire_0[107]);
  nand NAND2_256(keyinput_Wire_0[108], G642,G770);
  xor keyGate_0_108(G794, keyinput108, keyinput_Wire_0[108]);
  nand NAND2_257(G797,G645,G773);
  nand NAND2_258(G800,G648,G776);
  nand NAND2_259(keyinput_Wire_0[109], G651,G779);
  xor keyGate_0_109(KeyNOTWire_0[55], keyinput109, keyinput_Wire_0[109]);
  not KeyNOTGate_0_55(G803, KeyNOTWire_0[55]);
  nand NAND2_260(keyinput_Wire_0[110], G654,G782);
  xor keyGate_0_110(KeyNOTWire_0[56], keyinput110, keyinput_Wire_0[110]);
  not KeyNOTGate_0_56(G806, KeyNOTWire_0[56]);
  nand NAND2_261(keyinput_Wire_0[111], G657,G785);
  xnor keyGate_0_111(KeyNOTWire_0[57], keyinput111, keyinput_Wire_0[111]);
  not KeyNOTGate_0_57(G809, KeyNOTWire_0[57]);
  nand NAND2_262(G812,G660,G788);
  nand NAND2_263(G815,G663,G791);
  nand NAND2_264(G818,G642,G794);
  nand NAND2_265(G819,G770,G794);
  nand NAND2_266(G820,G645,G797);
  nand NAND2_267(G821,G773,G797);
  nand NAND2_268(keyinput_Wire_0[112], G648,G800);
  xor keyGate_0_112(G822, keyinput112, keyinput_Wire_0[112]);
  nand NAND2_269(G823,G776,G800);
  nand NAND2_270(keyinput_Wire_0[113], G651,G803);
  xnor keyGate_0_113(G824, keyinput113, keyinput_Wire_0[113]);
  nand NAND2_271(keyinput_Wire_0[114], G779,G803);
  xnor keyGate_0_114(G825, keyinput114, keyinput_Wire_0[114]);
  nand NAND2_272(G826,G654,G806);
  nand NAND2_273(G827,G782,G806);
  nand NAND2_274(keyinput_Wire_0[115], G657,G809);
  xnor keyGate_0_115(KeyNOTWire_0[58], keyinput115, keyinput_Wire_0[115]);
  not KeyNOTGate_0_58(G828, KeyNOTWire_0[58]);
  nand NAND2_275(keyinput_Wire_0[116], G785,G809);
  xor keyGate_0_116(KeyNOTWire_0[59], keyinput116, keyinput_Wire_0[116]);
  not KeyNOTGate_0_59(G829, KeyNOTWire_0[59]);
  nand NAND2_276(G830,G660,G812);
  nand NAND2_277(keyinput_Wire_0[117], G788,G812);
  xor keyGate_0_117(G831, keyinput117, keyinput_Wire_0[117]);
  nand NAND2_278(keyinput_Wire_0[118], G663,G815);
  xor keyGate_0_118(G832, keyinput118, keyinput_Wire_0[118]);
  nand NAND2_279(G833,G791,G815);
  nand NAND2_280(G834,G818,G819);
  nand NAND2_281(keyinput_Wire_0[119], G820,G821);
  xor keyGate_0_119(KeyNOTWire_0[60], keyinput119, keyinput_Wire_0[119]);
  not KeyNOTGate_0_60(G847, KeyNOTWire_0[60]);
  nand NAND2_282(keyinput_Wire_0[120], G822,G823);
  xnor keyGate_0_120(G860, keyinput120, keyinput_Wire_0[120]);
  nand NAND2_283(keyinput_Wire_0[121], G824,G825);
  xnor keyGate_0_121(G873, keyinput121, keyinput_Wire_0[121]);
  nand NAND2_284(G886,G828,G829);
  nand NAND2_285(keyinput_Wire_0[122], G832,G833);
  xnor keyGate_0_122(KeyNOTWire_0[61], keyinput122, keyinput_Wire_0[122]);
  not KeyNOTGate_0_61(G899, KeyNOTWire_0[61]);
  nand NAND2_286(G912,G830,G831);
  nand NAND2_287(G925,G826,G827);
  not NOT_0(G938,G834);
  not NOT_1(G939,G847);
  not NOT_2(G940,G860);
  not NOT_3(G941,G834);
  not NOT_4(G942,G847);
  not NOT_5(G943,G873);
  not NOT_6(G944,G834);
  not NOT_7(G945,G860);
  not NOT_8(G946,G873);
  not NOT_9(G947,G847);
  not NOT_10(G948,G860);
  not NOT_11(G949,G873);
  not NOT_12(G950,G886);
  not NOT_13(G951,G899);
  not NOT_14(G952,G886);
  not NOT_15(G953,G912);
  not NOT_16(G954,G925);
  not NOT_17(G955,G899);
  not NOT_18(G956,G925);
  not NOT_19(G957,G912);
  not NOT_20(G958,G925);
  not NOT_21(G959,G886);
  not NOT_22(G960,G912);
  not NOT_23(G961,G925);
  not NOT_24(G962,G886);
  not NOT_25(G963,G899);
  not NOT_26(G964,G925);
  not NOT_27(G965,G912);
  not NOT_28(G966,G899);
  not NOT_29(G967,G886);
  not NOT_30(G968,G912);
  not NOT_31(G969,G899);
  not NOT_32(G970,G847);
  not NOT_33(G971,G873);
  not NOT_34(G972,G847);
  not NOT_35(G973,G860);
  not NOT_36(G974,G834);
  not NOT_37(G975,G873);
  not NOT_38(G976,G834);
  not NOT_39(G977,G860);
  and AND4_0(G978,G938,G939,G940,G873);
  and AND4_1(G979,G941,G942,G860,G943);
  and AND4_2(G980,G944,G847,G945,G946);
  and AND4_3(G981,G834,G947,G948,G949);
  and AND4_4(G982,G958,G959,G960,G899);
  and AND4_5(G983,G961,G962,G912,G963);
  and AND4_6(G984,G964,G886,G965,G966);
  and AND4_7(G985,G925,G967,G968,G969);
  or OR4_0(G986,G978,G979,G980,G981);
  or OR4_1(G991,G982,G983,G984,G985);
  and AND5_0(G996,G925,G950,G912,G951,G986);
  and AND5_1(G1001,G925,G952,G953,G899,G986);
  and AND5_2(G1006,G954,G886,G912,G955,G986);
  and AND5_3(G1011,G956,G886,G957,G899,G986);
  and AND5_4(G1016,G834,G970,G860,G971,G991);
  and AND5_5(G1021,G834,G972,G973,G873,G991);
  and AND5_6(G1026,G974,G847,G860,G975,G991);
  and AND5_7(G1031,G976,G847,G977,G873,G991);
  and AND2_8(G1036,G834,G996);
  and AND2_9(G1039,G847,G996);
  and AND2_10(G1042,G860,G996);
  and AND2_11(G1045,G873,G996);
  and AND2_12(G1048,G834,G1001);
  and AND2_13(G1051,G847,G1001);
  and AND2_14(G1054,G860,G1001);
  and AND2_15(G1057,G873,G1001);
  and AND2_16(G1060,G834,G1006);
  and AND2_17(G1063,G847,G1006);
  and AND2_18(G1066,G860,G1006);
  and AND2_19(G1069,G873,G1006);
  and AND2_20(G1072,G834,G1011);
  and AND2_21(G1075,G847,G1011);
  and AND2_22(G1078,G860,G1011);
  and AND2_23(G1081,G873,G1011);
  and AND2_24(G1084,G925,G1016);
  and AND2_25(G1087,G886,G1016);
  and AND2_26(G1090,G912,G1016);
  and AND2_27(G1093,G899,G1016);
  and AND2_28(G1096,G925,G1021);
  and AND2_29(G1099,G886,G1021);
  and AND2_30(G1102,G912,G1021);
  and AND2_31(G1105,G899,G1021);
  and AND2_32(G1108,G925,G1026);
  and AND2_33(G1111,G886,G1026);
  and AND2_34(G1114,G912,G1026);
  and AND2_35(G1117,G899,G1026);
  and AND2_36(G1120,G925,G1031);
  and AND2_37(G1123,G886,G1031);
  and AND2_38(G1126,G912,G1031);
  and AND2_39(G1129,G899,G1031);
  nand NAND2_288(G1132,G1,G1036);
  nand NAND2_289(G1135,G2,G1039);
  nand NAND2_290(G1138,G3,G1042);
  nand NAND2_291(G1141,G4,G1045);
  nand NAND2_292(G1144,G5,G1048);
  nand NAND2_293(G1147,G6,G1051);
  nand NAND2_294(G1150,G7,G1054);
  nand NAND2_295(G1153,G8,G1057);
  nand NAND2_296(G1156,G9,G1060);
  nand NAND2_297(G1159,G10,G1063);
  nand NAND2_298(G1162,G11,G1066);
  nand NAND2_299(G1165,G12,G1069);
  nand NAND2_300(G1168,G13,G1072);
  nand NAND2_301(G1171,G14,G1075);
  nand NAND2_302(G1174,G15,G1078);
  nand NAND2_303(G1177,G16,G1081);
  nand NAND2_304(G1180,G17,G1084);
  nand NAND2_305(G1183,G18,G1087);
  nand NAND2_306(G1186,G19,G1090);
  nand NAND2_307(keyinput_Wire_0[123], G20,G1093);
  xor keyGate_0_123(G1189, keyinput123, keyinput_Wire_0[123]);
  nand NAND2_308(G1192,G21,G1096);
  nand NAND2_309(G1195,G22,G1099);
  nand NAND2_310(G1198,G23,G1102);
  nand NAND2_311(G1201,G24,G1105);
  nand NAND2_312(G1204,G25,G1108);
  nand NAND2_313(G1207,G26,G1111);
  nand NAND2_314(G1210,G27,G1114);
  nand NAND2_315(G1213,G28,G1117);
  nand NAND2_316(G1216,G29,G1120);
  nand NAND2_317(G1219,G30,G1123);
  nand NAND2_318(G1222,G31,G1126);
  nand NAND2_319(G1225,G32,G1129);
  nand NAND2_320(G1228,G1,G1132);
  nand NAND2_321(G1229,G1036,G1132);
  nand NAND2_322(G1230,G2,G1135);
  nand NAND2_323(G1231,G1039,G1135);
  nand NAND2_324(G1232,G3,G1138);
  nand NAND2_325(G1233,G1042,G1138);
  nand NAND2_326(G1234,G4,G1141);
  nand NAND2_327(G1235,G1045,G1141);
  nand NAND2_328(G1236,G5,G1144);
  nand NAND2_329(keyinput_Wire_0[124], G1048,G1144);
  xor keyGate_0_124(KeyNOTWire_0[62], keyinput124, keyinput_Wire_0[124]);
  not KeyNOTGate_0_62(G1237, KeyNOTWire_0[62]);
  nand NAND2_330(G1238,G6,G1147);
  nand NAND2_331(G1239,G1051,G1147);
  nand NAND2_332(G1240,G7,G1150);
  nand NAND2_333(G1241,G1054,G1150);
  nand NAND2_334(G1242,G8,G1153);
  nand NAND2_335(G1243,G1057,G1153);
  nand NAND2_336(G1244,G9,G1156);
  nand NAND2_337(G1245,G1060,G1156);
  nand NAND2_338(keyinput_Wire_0[125], G10,G1159);
  xor keyGate_0_125(KeyNOTWire_0[63], keyinput125, keyinput_Wire_0[125]);
  not KeyNOTGate_0_63(G1246, KeyNOTWire_0[63]);
  nand NAND2_339(G1247,G1063,G1159);
  nand NAND2_340(keyinput_Wire_0[126], G11,G1162);
  xor keyGate_0_126(KeyNOTWire_0[64], keyinput126, keyinput_Wire_0[126]);
  not KeyNOTGate_0_64(G1248, KeyNOTWire_0[64]);
  nand NAND2_341(G1249,G1066,G1162);
  nand NAND2_342(G1250,G12,G1165);
  nand NAND2_343(G1251,G1069,G1165);
  nand NAND2_344(keyinput_Wire_0[127], G13,G1168);
  xnor keyGate_0_127(G1252, keyinput127, keyinput_Wire_0[127]);
  nand NAND2_345(G1253,G1072,G1168);
  nand NAND2_346(G1254,G14,G1171);
  nand NAND2_347(G1255,G1075,G1171);
  nand NAND2_348(G1256,G15,G1174);
  nand NAND2_349(G1257,G1078,G1174);
  nand NAND2_350(G1258,G16,G1177);
  nand NAND2_351(G1259,G1081,G1177);
  nand NAND2_352(G1260,G17,G1180);
  nand NAND2_353(G1261,G1084,G1180);
  nand NAND2_354(G1262,G18,G1183);
  nand NAND2_355(G1263,G1087,G1183);
  nand NAND2_356(G1264,G19,G1186);
  nand NAND2_357(G1265,G1090,G1186);
  nand NAND2_358(G1266,G20,G1189);
  nand NAND2_359(G1267,G1093,G1189);
  nand NAND2_360(G1268,G21,G1192);
  nand NAND2_361(G1269,G1096,G1192);
  nand NAND2_362(G1270,G22,G1195);
  nand NAND2_363(G1271,G1099,G1195);
  nand NAND2_364(G1272,G23,G1198);
  nand NAND2_365(G1273,G1102,G1198);
  nand NAND2_366(G1274,G24,G1201);
  nand NAND2_367(G1275,G1105,G1201);
  nand NAND2_368(G1276,G25,G1204);
  nand NAND2_369(G1277,G1108,G1204);
  nand NAND2_370(G1278,G26,G1207);
  nand NAND2_371(G1279,G1111,G1207);
  nand NAND2_372(G1280,G27,G1210);
  nand NAND2_373(G1281,G1114,G1210);
  nand NAND2_374(G1282,G28,G1213);
  nand NAND2_375(G1283,G1117,G1213);
  nand NAND2_376(G1284,G29,G1216);
  nand NAND2_377(G1285,G1120,G1216);
  nand NAND2_378(G1286,G30,G1219);
  nand NAND2_379(G1287,G1123,G1219);
  nand NAND2_380(G1288,G31,G1222);
  nand NAND2_381(G1289,G1126,G1222);
  nand NAND2_382(G1290,G32,G1225);
  nand NAND2_383(G1291,G1129,G1225);
  nand NAND2_384(G1292,G1228,G1229);
  nand NAND2_385(G1293,G1230,G1231);
  nand NAND2_386(G1294,G1232,G1233);
  nand NAND2_387(G1295,G1234,G1235);
  nand NAND2_388(G1296,G1236,G1237);
  nand NAND2_389(G1297,G1238,G1239);
  nand NAND2_390(G1298,G1240,G1241);
  nand NAND2_391(G1299,G1242,G1243);
  nand NAND2_392(G1300,G1244,G1245);
  nand NAND2_393(G1301,G1246,G1247);
  nand NAND2_394(G1302,G1248,G1249);
  nand NAND2_395(G1303,G1250,G1251);
  nand NAND2_396(G1304,G1252,G1253);
  nand NAND2_397(G1305,G1254,G1255);
  nand NAND2_398(G1306,G1256,G1257);
  nand NAND2_399(G1307,G1258,G1259);
  nand NAND2_400(G1308,G1260,G1261);
  nand NAND2_401(G1309,G1262,G1263);
  nand NAND2_402(G1310,G1264,G1265);
  nand NAND2_403(G1311,G1266,G1267);
  nand NAND2_404(G1312,G1268,G1269);
  nand NAND2_405(G1313,G1270,G1271);
  nand NAND2_406(G1314,G1272,G1273);
  nand NAND2_407(G1315,G1274,G1275);
  nand NAND2_408(G1316,G1276,G1277);
  nand NAND2_409(G1317,G1278,G1279);
  nand NAND2_410(G1318,G1280,G1281);
  nand NAND2_411(G1319,G1282,G1283);
  nand NAND2_412(G1320,G1284,G1285);
  nand NAND2_413(G1321,G1286,G1287);
  nand NAND2_414(G1322,G1288,G1289);
  nand NAND2_415(G1323,G1290,G1291);
  not NOT_40(G1324,G1292);
  not NOT_41(G1325,G1293);
  not NOT_42(G1326,G1294);
  not NOT_43(G1327,G1295);
  not NOT_44(G1328,G1296);
  not NOT_45(G1329,G1297);
  not NOT_46(G1330,G1298);
  not NOT_47(KeyWire_0_1,G1299);
  xor flip_it (G1331, KeyWire_0_1, KeyWire_0_2 );
  not NOT_48(G1332,G1300);
  not NOT_49(G1333,G1301);
  not NOT_50(G1334,G1302);
  not NOT_51(G1335,G1303);
  not NOT_52(G1336,G1304);
  not NOT_53(G1337,G1305);
  not NOT_54(G1338,G1306);
  not NOT_55(G1339,G1307);
  not NOT_56(G1340,G1308);
  not NOT_57(G1341,G1309);
  not NOT_58(G1342,G1310);
  not NOT_59(G1343,G1311);
  not NOT_60(G1344,G1312);
  not NOT_61(G1345,G1313);
  not NOT_62(G1346,G1314);
  not NOT_63(G1347,G1315);
  not NOT_64(G1348,G1316);
  not NOT_65(G1349,G1317);
  not NOT_66(G1350,G1318);
  not NOT_67(G1351,G1319);
  not NOT_68(G1352,G1320);
  not NOT_69(G1353,G1321);
  not NOT_70(G1354,G1322);
  not NOT_71(G1355,G1323);

AntiSAT some_name( KeyWire_0_2, G36, G32, G18, G21, G25, G26, G27, G24, G20, G23, G35, G8, G30, G31, G10, G1, G7, G6, G14, G40, G4, G34, G12, G16, G17, G19, G41, G33, G11, G22, G29, G15, G3, G37, G9, G13, G2, G38, G5, G28, G39, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
       keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
       keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
       keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
       keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
       keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
       keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
       keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
       keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
       keyinput250);

endmodule


/*************************************************************************/

module AntiSAT (KeyWire_0_2, G36, G32, G18, G21, G25, G26, G27, G24, G20, G23, G35, G8, G30, G31, G10, G1, G7, G6, G14, G40, G4, G34, G12, G16, G17, G19, G41, G33, G11, G22, G29, G15, G3, G37, G9, G13, G2, G38, G5, G28, G39, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, keyinput208, keyinput209 ,
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
        keyinput250);

  input keyinput210, keyinput211, keyinput212, keyinput213, keyinput214;
  input keyinput215, keyinput216, keyinput217, keyinput218, keyinput219;
  input keyinput220, keyinput221, keyinput222, keyinput223, keyinput224;
  input keyinput225, keyinput226, keyinput227, keyinput228, keyinput229;
  input keyinput230, keyinput231, keyinput232, keyinput233, keyinput234;
  input keyinput235, keyinput236, keyinput237, keyinput238, keyinput239;
  input keyinput240, keyinput241, keyinput242, keyinput243, keyinput244;
  input keyinput245, keyinput246, keyinput247, keyinput248, keyinput249;
  input keyinput250;

  wire [0:40] keyNTin_Wire_1;
  wire [0:22] KeyNOTWire_1;

  input G36, G32, G18, G21, G25, G26, G27, G24, G20, G23, G35, G8, G30, G31, G10, G1, G7, G6, G14, G40, G4, G34, G12, G16, G17, G19, G41, G33, G11, G22, G29, G15, G3, G37, G9, G13, G2, G38, G5, G28, G39;
  input keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, keyinput208, keyinput209;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83 ;

  xnor KeyGate0 (keyNTin_Wire_1[0], G36, keyinput128);
  xor keyNTinGate_1_0(KeyNOTWire_1[0], keyinput210, keyNTin_Wire_1[0]);
  not KeyNOTGate_1_0(newWire_0, KeyNOTWire_1[0]);
  xor  KeyGate1 (newWire_1, G32, keyinput129);
  xnor KeyGate2 (newWire_2, G18, keyinput130);
  xor  KeyGate3 (newWire_3, G21, keyinput131);
  xnor KeyGate4 (newWire_4, G25, keyinput132);
  xnor KeyGate5 (keyNTin_Wire_1[1], G26, keyinput133);
  xnor keyNTinGate_1_1(KeyNOTWire_1[1], keyinput211, keyNTin_Wire_1[1]);
  not KeyNOTGate_1_1(newWire_5, KeyNOTWire_1[1]);
  xor  KeyGate6 (newWire_6, G27, keyinput134);
  xor  KeyGate7 (keyNTin_Wire_1[2], G24, keyinput135);
  xnor keyNTinGate_1_2(KeyNOTWire_1[2], keyinput212, keyNTin_Wire_1[2]);
  not KeyNOTGate_1_2(newWire_7, KeyNOTWire_1[2]);
  xnor KeyGate8 (newWire_8, G20, keyinput136);
  xnor KeyGate9 (keyNTin_Wire_1[3], G23, keyinput137);
  xor keyNTinGate_1_3(KeyNOTWire_1[3], keyinput213, keyNTin_Wire_1[3]);
  not KeyNOTGate_1_3(newWire_9, KeyNOTWire_1[3]);
  xnor KeyGate10 (keyNTin_Wire_1[4], G35, keyinput138);
  xnor keyNTinGate_1_4(newWire_10, keyinput214, keyNTin_Wire_1[4]);
  xnor KeyGate11 (keyNTin_Wire_1[5], G8, keyinput139);
  xnor keyNTinGate_1_5(newWire_11, keyinput215, keyNTin_Wire_1[5]);
  xor  KeyGate12 (keyNTin_Wire_1[6], G30, keyinput140);
  xor keyNTinGate_1_6(KeyNOTWire_1[4], keyinput216, keyNTin_Wire_1[6]);
  not KeyNOTGate_1_4(newWire_12, KeyNOTWire_1[4]);
  xor  KeyGate13 (keyNTin_Wire_1[7], G31, keyinput141);
  xor keyNTinGate_1_7(KeyNOTWire_1[5], keyinput217, keyNTin_Wire_1[7]);
  not KeyNOTGate_1_5(newWire_13, KeyNOTWire_1[5]);
  xor  KeyGate14 (newWire_14, G10, keyinput142);
  xnor KeyGate15 (newWire_15, G1, keyinput143);
  xnor KeyGate16 (newWire_16, G7, keyinput144);
  xor  KeyGate17 (keyNTin_Wire_1[8], G6, keyinput145);
  xnor keyNTinGate_1_8(KeyNOTWire_1[6], keyinput218, keyNTin_Wire_1[8]);
  not KeyNOTGate_1_6(newWire_17, KeyNOTWire_1[6]);
  xor  KeyGate18 (newWire_18, G14, keyinput146);
  xnor KeyGate19 (newWire_19, G40, keyinput147);
  xnor KeyGate20 (newWire_20, G4, keyinput148);
  xnor KeyGate21 (newWire_21, G34, keyinput149);
  xnor KeyGate22 (newWire_22, G12, keyinput150);
  xnor KeyGate23 (newWire_23, G16, keyinput151);
  xor  KeyGate24 (keyNTin_Wire_1[9], G17, keyinput152);
  xnor keyNTinGate_1_9(newWire_24, keyinput219, keyNTin_Wire_1[9]);
  xnor KeyGate25 (newWire_25, G19, keyinput153);
  xor  KeyGate26 (keyNTin_Wire_1[10], G41, keyinput154);
  xnor keyNTinGate_1_10(newWire_26, keyinput220, keyNTin_Wire_1[10]);
  xnor KeyGate27 (newWire_27, G33, keyinput155);
  xnor KeyGate28 (newWire_28, G11, keyinput156);
  xor  KeyGate29 (keyNTin_Wire_1[11], G22, keyinput157);
  xnor keyNTinGate_1_11(newWire_29, keyinput221, keyNTin_Wire_1[11]);
  xor  KeyGate30 (keyNTin_Wire_1[12], G29, keyinput158);
  xor keyNTinGate_1_12(newWire_30, keyinput222, keyNTin_Wire_1[12]);
  xnor KeyGate31 (newWire_31, G15, keyinput159);
  xnor KeyGate32 (newWire_32, G3, keyinput160);
  xnor KeyGate33 (newWire_33, G37, keyinput161);
  xor  KeyGate34 (newWire_34, G9, keyinput162);
  xnor KeyGate35 (keyNTin_Wire_1[13], G13, keyinput163);
  xor keyNTinGate_1_13(newWire_35, keyinput223, keyNTin_Wire_1[13]);
  xor  KeyGate36 (newWire_36, G2, keyinput164);
  xnor KeyGate37 (newWire_37, G38, keyinput165);
  xnor KeyGate38 (keyNTin_Wire_1[14], G5, keyinput166);
  xnor keyNTinGate_1_14(KeyNOTWire_1[7], keyinput224, keyNTin_Wire_1[14]);
  not KeyNOTGate_1_7(newWire_38, KeyNOTWire_1[7]);
  xor  KeyGate39 (newWire_39, G28, keyinput167);
  xnor KeyGate40 (newWire_40, G39, keyinput168);
  xnor KeyGate41 (newWire_41, G36, keyinput169);
  xnor KeyGate42 (keyNTin_Wire_1[15], G32, keyinput170);
  xor keyNTinGate_1_15(KeyNOTWire_1[8], keyinput225, keyNTin_Wire_1[15]);
  not KeyNOTGate_1_8(newWire_42, KeyNOTWire_1[8]);
  xor  KeyGate43 (keyNTin_Wire_1[16], G18, keyinput171);
  xnor keyNTinGate_1_16(KeyNOTWire_1[9], keyinput226, keyNTin_Wire_1[16]);
  not KeyNOTGate_1_9(newWire_43, KeyNOTWire_1[9]);
  xnor KeyGate44 (keyNTin_Wire_1[17], G21, keyinput172);
  xor keyNTinGate_1_17(KeyNOTWire_1[10], keyinput227, keyNTin_Wire_1[17]);
  not KeyNOTGate_1_10(newWire_44, KeyNOTWire_1[10]);
  xor  KeyGate45 (keyNTin_Wire_1[18], G25, keyinput173);
  xor keyNTinGate_1_18(KeyNOTWire_1[11], keyinput228, keyNTin_Wire_1[18]);
  not KeyNOTGate_1_11(newWire_45, KeyNOTWire_1[11]);
  xor  KeyGate46 (newWire_46, G26, keyinput174);
  xnor KeyGate47 (keyNTin_Wire_1[19], G27, keyinput175);
  xnor keyNTinGate_1_19(newWire_47, keyinput229, keyNTin_Wire_1[19]);
  xnor KeyGate48 (newWire_48, G24, keyinput176);
  xnor KeyGate49 (newWire_49, G20, keyinput177);
  xnor KeyGate50 (newWire_50, G23, keyinput178);
  xnor KeyGate51 (keyNTin_Wire_1[20], G35, keyinput179);
  xnor keyNTinGate_1_20(KeyNOTWire_1[12], keyinput230, keyNTin_Wire_1[20]);
  not KeyNOTGate_1_12(newWire_51, KeyNOTWire_1[12]);
  xor  KeyGate52 (keyNTin_Wire_1[21], G8, keyinput180);
  xor keyNTinGate_1_21(KeyNOTWire_1[13], keyinput231, keyNTin_Wire_1[21]);
  not KeyNOTGate_1_13(newWire_52, KeyNOTWire_1[13]);
  xnor KeyGate53 (newWire_53, G30, keyinput181);
  xnor KeyGate54 (newWire_54, G31, keyinput182);
  xnor KeyGate55 (keyNTin_Wire_1[22], G10, keyinput183);
  xor keyNTinGate_1_22(KeyNOTWire_1[14], keyinput232, keyNTin_Wire_1[22]);
  not KeyNOTGate_1_14(newWire_55, KeyNOTWire_1[14]);
  xnor KeyGate56 (keyNTin_Wire_1[23], G1, keyinput184);
  xor keyNTinGate_1_23(newWire_56, keyinput233, keyNTin_Wire_1[23]);
  xor  KeyGate57 (keyNTin_Wire_1[24], G7, keyinput185);
  xor keyNTinGate_1_24(KeyNOTWire_1[15], keyinput234, keyNTin_Wire_1[24]);
  not KeyNOTGate_1_15(newWire_57, KeyNOTWire_1[15]);
  xnor KeyGate58 (keyNTin_Wire_1[25], G6, keyinput186);
  xor keyNTinGate_1_25(newWire_58, keyinput235, keyNTin_Wire_1[25]);
  xor  KeyGate59 (keyNTin_Wire_1[26], G14, keyinput187);
  xnor keyNTinGate_1_26(KeyNOTWire_1[16], keyinput236, keyNTin_Wire_1[26]);
  not KeyNOTGate_1_16(newWire_59, KeyNOTWire_1[16]);
  xor  KeyGate60 (keyNTin_Wire_1[27], G40, keyinput188);
  xnor keyNTinGate_1_27(KeyNOTWire_1[17], keyinput237, keyNTin_Wire_1[27]);
  not KeyNOTGate_1_17(newWire_60, KeyNOTWire_1[17]);
  xor  KeyGate61 (keyNTin_Wire_1[28], G4, keyinput189);
  xnor keyNTinGate_1_28(newWire_61, keyinput238, keyNTin_Wire_1[28]);
  xnor KeyGate62 (newWire_62, G34, keyinput190);
  xor  KeyGate63 (keyNTin_Wire_1[29], G12, keyinput191);
  xor keyNTinGate_1_29(newWire_63, keyinput239, keyNTin_Wire_1[29]);
  xnor KeyGate64 (keyNTin_Wire_1[30], G16, keyinput192);
  xnor keyNTinGate_1_30(newWire_64, keyinput240, keyNTin_Wire_1[30]);
  xor  KeyGate65 (keyNTin_Wire_1[31], G17, keyinput193);
  xor keyNTinGate_1_31(KeyNOTWire_1[18], keyinput241, keyNTin_Wire_1[31]);
  not KeyNOTGate_1_18(newWire_65, KeyNOTWire_1[18]);
  xor  KeyGate66 (keyNTin_Wire_1[32], G19, keyinput194);
  xnor keyNTinGate_1_32(KeyNOTWire_1[19], keyinput242, keyNTin_Wire_1[32]);
  not KeyNOTGate_1_19(newWire_66, KeyNOTWire_1[19]);
  xor  KeyGate67 (keyNTin_Wire_1[33], G41, keyinput195);
  xnor keyNTinGate_1_33(newWire_67, keyinput243, keyNTin_Wire_1[33]);
  xnor KeyGate68 (newWire_68, G33, keyinput196);
  xnor KeyGate69 (keyNTin_Wire_1[34], G11, keyinput197);
  xnor keyNTinGate_1_34(KeyNOTWire_1[20], keyinput244, keyNTin_Wire_1[34]);
  not KeyNOTGate_1_20(newWire_69, KeyNOTWire_1[20]);
  xnor KeyGate70 (keyNTin_Wire_1[35], G22, keyinput198);
  xor keyNTinGate_1_35(newWire_70, keyinput245, keyNTin_Wire_1[35]);
  xnor KeyGate71 (keyNTin_Wire_1[36], G29, keyinput199);
  xor keyNTinGate_1_36(newWire_71, keyinput246, keyNTin_Wire_1[36]);
  xor  KeyGate72 (keyNTin_Wire_1[37], G15, keyinput200);
  xnor keyNTinGate_1_37(newWire_72, keyinput247, keyNTin_Wire_1[37]);
  xor  KeyGate73 (newWire_73, G3, keyinput201);
  xnor KeyGate74 (newWire_74, G37, keyinput202);
  xnor KeyGate75 (newWire_75, G9, keyinput203);
  xor  KeyGate76 (keyNTin_Wire_1[38], G13, keyinput204);
  xor keyNTinGate_1_38(newWire_76, keyinput248, keyNTin_Wire_1[38]);
  xnor KeyGate77 (newWire_77, G2, keyinput205);
  xor  KeyGate78 (keyNTin_Wire_1[39], G38, keyinput206);
  xnor keyNTinGate_1_39(KeyNOTWire_1[21], keyinput249, keyNTin_Wire_1[39]);
  not KeyNOTGate_1_21(newWire_78, KeyNOTWire_1[21]);
  xor  KeyGate79 (newWire_79, G5, keyinput207);
  xor  KeyGate80 (newWire_80, G28, keyinput208);
  xnor KeyGate81 (newWire_81, G39, keyinput209);
  and some_function (newWire_82, newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40 );
  nand compl_function (newWire_83, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81);
  and finalAND (keyNTin_Wire_1[40], newWire_82, newWire_83);
  xor keyNTinGate_1_40(KeyNOTWire_1[22], keyinput250, keyNTin_Wire_1[40]);
  not KeyNOTGate_1_22(KeyWire_0_2, KeyNOTWire_1[22]);

endmodule /* AntiSAT */
