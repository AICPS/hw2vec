`timescale 1ns / 1ps
// Verilog
// c499
// Ninputs 41
// Noutputs 32
// NtotalGates 202
// XOR2 104
// AND2 40
// NOT1 40
// AND4 8
// OR4 2
// AND5 8

module top (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
                  N753,N754,N755,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
                  keyinput60, keyinput61, keyinput62, keyinput63,
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
        keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
        keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
        keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
        keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
        keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
        keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
        keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
                  keyinput144, keyinput145,
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150,
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155,
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160,
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165,
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170,
        keyinput171, keyinput172, keyinput173, keyinput174, keyinput175,
        keyinput176, keyinput177, keyinput178, keyinput179, keyinput180,
        keyinput181, keyinput182, keyinput183, keyinput184, keyinput185,
        keyinput186);

  input keyinput146, keyinput147, keyinput148, keyinput149, keyinput150;
  input keyinput151, keyinput152, keyinput153, keyinput154, keyinput155;
  input keyinput156, keyinput157, keyinput158, keyinput159, keyinput160;
  input keyinput161, keyinput162, keyinput163, keyinput164, keyinput165;
  input keyinput166, keyinput167, keyinput168, keyinput169, keyinput170;
  input keyinput171, keyinput172, keyinput173, keyinput174, keyinput175;
  input keyinput176, keyinput177, keyinput178, keyinput179, keyinput180;
  input keyinput181, keyinput182, keyinput183, keyinput184, keyinput185;
  input keyinput186;


  input keyinput64, keyinput65, keyinput66, keyinput67, keyinput68;
  input keyinput69, keyinput70, keyinput71, keyinput72, keyinput73;
  input keyinput74, keyinput75, keyinput76, keyinput77, keyinput78;
  input keyinput79, keyinput80, keyinput81, keyinput82, keyinput83;
  input keyinput84, keyinput85, keyinput86, keyinput87, keyinput88;
  input keyinput89, keyinput90, keyinput91, keyinput92, keyinput93;
  input keyinput94, keyinput95, keyinput96, keyinput97, keyinput98;
  input keyinput99, keyinput100, keyinput101, keyinput102, keyinput103;
  input keyinput104, keyinput105, keyinput106, keyinput107, keyinput108;
  input keyinput109, keyinput110, keyinput111, keyinput112, keyinput113;
  input keyinput114, keyinput115, keyinput116, keyinput117, keyinput118;
  input keyinput119, keyinput120, keyinput121, keyinput122, keyinput123;
  input keyinput124, keyinput125, keyinput126, keyinput127, keyinput128;
  input keyinput129, keyinput130, keyinput131, keyinput132, keyinput133;
  input keyinput134, keyinput135, keyinput136, keyinput137, keyinput138;
  input keyinput139, keyinput140, keyinput141, keyinput142, keyinput143;
  input keyinput144, keyinput145;

  wire KeyWire_0_1 , KeyWire_0_2;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31, keyinput32, keyinput33, keyinput34;
  input keyinput35, keyinput36, keyinput37, keyinput38, keyinput39;
  input keyinput40, keyinput41, keyinput42, keyinput43, keyinput44;
  input keyinput45, keyinput46, keyinput47, keyinput48, keyinput49;
  input keyinput50, keyinput51, keyinput52, keyinput53, keyinput54;
  input keyinput55, keyinput56, keyinput57, keyinput58, keyinput59;
  input keyinput60, keyinput61, keyinput62, keyinput63;

  wire [0:63] keyinput_Wire_0;
  wire [0:32] KeyNOTWire_0;

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;

output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723;

  xor XOR2_1 (keyinput_Wire_0[0], N1, N5);
  xor keyGate_0_0(KeyNOTWire_0[0], keyinput0, keyinput_Wire_0[0]);
  not KeyNOTGate_0_0(N250, KeyNOTWire_0[0]);
xor XOR2_2 (N251, N9, N13);
  xor XOR2_3 (keyinput_Wire_0[1], N17, N21);
  xnor keyGate_0_1(N252, keyinput1, keyinput_Wire_0[1]);
  xor XOR2_4 (keyinput_Wire_0[2], N25, N29);
  xor keyGate_0_2(KeyNOTWire_0[1], keyinput2, keyinput_Wire_0[2]);
  not KeyNOTGate_0_1(N253, KeyNOTWire_0[1]);
xor XOR2_5 (N254, N33, N37);
  xor XOR2_6 (keyinput_Wire_0[3], N41, N45);
  xnor keyGate_0_3(N255, keyinput3, keyinput_Wire_0[3]);
  xor XOR2_7 (keyinput_Wire_0[4], N49, N53);
  xnor keyGate_0_4(KeyNOTWire_0[2], keyinput4, keyinput_Wire_0[4]);
  not KeyNOTGate_0_2(N256, KeyNOTWire_0[2]);
  xor XOR2_8 (keyinput_Wire_0[5], N57, N61);
  xnor keyGate_0_5(N257, keyinput5, keyinput_Wire_0[5]);
xor XOR2_9 (N258, N65, N69);
  xor XOR2_10 (keyinput_Wire_0[6], N73, N77);
  xor keyGate_0_6(KeyNOTWire_0[3], keyinput6, keyinput_Wire_0[6]);
  not KeyNOTGate_0_3(N259, KeyNOTWire_0[3]);
  xor XOR2_11 (keyinput_Wire_0[7], N81, N85);
  xor keyGate_0_7(KeyNOTWire_0[4], keyinput7, keyinput_Wire_0[7]);
  not KeyNOTGate_0_4(N260, KeyNOTWire_0[4]);
  xor XOR2_12 (keyinput_Wire_0[8], N89, N93);
  xor keyGate_0_8(N261, keyinput8, keyinput_Wire_0[8]);
  xor XOR2_13 (keyinput_Wire_0[9], N97, N101);
  xnor keyGate_0_9(KeyNOTWire_0[5], keyinput9, keyinput_Wire_0[9]);
  not KeyNOTGate_0_5(N262, KeyNOTWire_0[5]);
  xor XOR2_14 (keyinput_Wire_0[10], N105, N109);
  xor keyGate_0_10(KeyNOTWire_0[6], keyinput10, keyinput_Wire_0[10]);
  not KeyNOTGate_0_6(N263, KeyNOTWire_0[6]);
xor XOR2_15 (N264, N113, N117);
xor XOR2_16 (N265, N121, N125);
  and AND2_17 (keyinput_Wire_0[11], N129, N137);
  xor keyGate_0_11(N266, keyinput11, keyinput_Wire_0[11]);
  and AND2_18 (keyinput_Wire_0[12], N130, N137);
  xnor keyGate_0_12(KeyNOTWire_0[7], keyinput12, keyinput_Wire_0[12]);
  not KeyNOTGate_0_7(N267, KeyNOTWire_0[7]);
  and AND2_19 (keyinput_Wire_0[13], N131, N137);
  xnor keyGate_0_13(N268, keyinput13, keyinput_Wire_0[13]);
and AND2_20 (N269, N132, N137);
  and AND2_21 (keyinput_Wire_0[14], N133, N137);
  xor keyGate_0_14(KeyNOTWire_0[8], keyinput14, keyinput_Wire_0[14]);
  not KeyNOTGate_0_8(N270, KeyNOTWire_0[8]);
  and AND2_22 (keyinput_Wire_0[15], N134, N137);
  xor keyGate_0_15(KeyNOTWire_0[9], keyinput15, keyinput_Wire_0[15]);
  not KeyNOTGate_0_9(N271, KeyNOTWire_0[9]);
  and AND2_23 (keyinput_Wire_0[16], N135, N137);
  xnor keyGate_0_16(N272, keyinput16, keyinput_Wire_0[16]);
  and AND2_24 (keyinput_Wire_0[17], N136, N137);
  xnor keyGate_0_17(N273, keyinput17, keyinput_Wire_0[17]);
  xor XOR2_25 (keyinput_Wire_0[18], N1, N17);
  xnor keyGate_0_18(N274, keyinput18, keyinput_Wire_0[18]);
xor XOR2_26 (N275, N33, N49);
xor XOR2_27 (N276, N5, N21);
  xor XOR2_28 (keyinput_Wire_0[19], N37, N53);
  xnor keyGate_0_19(N277, keyinput19, keyinput_Wire_0[19]);
  xor XOR2_29 (keyinput_Wire_0[20], N9, N25);
  xnor keyGate_0_20(KeyNOTWire_0[10], keyinput20, keyinput_Wire_0[20]);
  not KeyNOTGate_0_10(N278, KeyNOTWire_0[10]);
xor XOR2_30 (N279, N41, N57);
  xor XOR2_31 (keyinput_Wire_0[21], N13, N29);
  xnor keyGate_0_21(KeyNOTWire_0[11], keyinput21, keyinput_Wire_0[21]);
  not KeyNOTGate_0_11(N280, KeyNOTWire_0[11]);
  xor XOR2_32 (keyinput_Wire_0[22], N45, N61);
  xor keyGate_0_22(KeyNOTWire_0[12], keyinput22, keyinput_Wire_0[22]);
  not KeyNOTGate_0_12(N281, KeyNOTWire_0[12]);
  xor XOR2_33 (keyinput_Wire_0[23], N65, N81);
  xor keyGate_0_23(N282, keyinput23, keyinput_Wire_0[23]);
  xor XOR2_34 (keyinput_Wire_0[24], N97, N113);
  xnor keyGate_0_24(KeyNOTWire_0[13], keyinput24, keyinput_Wire_0[24]);
  not KeyNOTGate_0_13(N283, KeyNOTWire_0[13]);
  xor XOR2_35 (keyinput_Wire_0[25], N69, N85);
  xor keyGate_0_25(KeyNOTWire_0[14], keyinput25, keyinput_Wire_0[25]);
  not KeyNOTGate_0_14(N284, KeyNOTWire_0[14]);
  xor XOR2_36 (keyinput_Wire_0[26], N101, N117);
  xnor keyGate_0_26(N285, keyinput26, keyinput_Wire_0[26]);
  xor XOR2_37 (keyinput_Wire_0[27], N73, N89);
  xnor keyGate_0_27(N286, keyinput27, keyinput_Wire_0[27]);
  xor XOR2_38 (keyinput_Wire_0[28], N105, N121);
  xnor keyGate_0_28(KeyNOTWire_0[15], keyinput28, keyinput_Wire_0[28]);
  not KeyNOTGate_0_15(N287, KeyNOTWire_0[15]);
  xor XOR2_39 (keyinput_Wire_0[29], N77, N93);
  xnor keyGate_0_29(KeyNOTWire_0[16], keyinput29, keyinput_Wire_0[29]);
  not KeyNOTGate_0_16(N288, KeyNOTWire_0[16]);
  xor XOR2_40 (keyinput_Wire_0[30], N109, N125);
  xnor keyGate_0_30(N289, keyinput30, keyinput_Wire_0[30]);
xor XOR2_41 (N290, N250, N251);
  xor XOR2_42 (keyinput_Wire_0[31], N252, N253);
  xor keyGate_0_31(KeyNOTWire_0[17], keyinput31, keyinput_Wire_0[31]);
  not KeyNOTGate_0_17(N293, KeyNOTWire_0[17]);
  xor XOR2_43 (keyinput_Wire_0[32], N254, N255);
  xor keyGate_0_32(N296, keyinput32, keyinput_Wire_0[32]);
  xor XOR2_44 (keyinput_Wire_0[33], N256, N257);
  xor keyGate_0_33(N299, keyinput33, keyinput_Wire_0[33]);
xor XOR2_45 (N302, N258, N259);
  xor XOR2_46 (keyinput_Wire_0[34], N260, N261);
  xnor keyGate_0_34(KeyNOTWire_0[18], keyinput34, keyinput_Wire_0[34]);
  not KeyNOTGate_0_18(N305, KeyNOTWire_0[18]);
  xor XOR2_47 (keyinput_Wire_0[35], N262, N263);
  xor keyGate_0_35(N308, keyinput35, keyinput_Wire_0[35]);
xor XOR2_48 (N311, N264, N265);
  xor XOR2_49 (keyinput_Wire_0[36], N274, N275);
  xor keyGate_0_36(N314, keyinput36, keyinput_Wire_0[36]);
  xor XOR2_50 (keyinput_Wire_0[37], N276, N277);
  xnor keyGate_0_37(KeyNOTWire_0[19], keyinput37, keyinput_Wire_0[37]);
  not KeyNOTGate_0_19(N315, KeyNOTWire_0[19]);
  xor XOR2_51 (keyinput_Wire_0[38], N278, N279);
  xor keyGate_0_38(KeyNOTWire_0[20], keyinput38, keyinput_Wire_0[38]);
  not KeyNOTGate_0_20(N316, KeyNOTWire_0[20]);
  xor XOR2_52 (keyinput_Wire_0[39], N280, N281);
  xor keyGate_0_39(KeyNOTWire_0[21], keyinput39, keyinput_Wire_0[39]);
  not KeyNOTGate_0_21(N317, KeyNOTWire_0[21]);
  xor XOR2_53 (keyinput_Wire_0[40], N282, N283);
  xnor keyGate_0_40(KeyNOTWire_0[22], keyinput40, keyinput_Wire_0[40]);
  not KeyNOTGate_0_22(N318, KeyNOTWire_0[22]);
  xor XOR2_54 (keyinput_Wire_0[41], N284, N285);
  xnor keyGate_0_41(N319, keyinput41, keyinput_Wire_0[41]);
  xor XOR2_55 (keyinput_Wire_0[42], N286, N287);
  xnor keyGate_0_42(KeyNOTWire_0[23], keyinput42, keyinput_Wire_0[42]);
  not KeyNOTGate_0_23(N320, KeyNOTWire_0[23]);
  xor XOR2_56 (keyinput_Wire_0[43], N288, N289);
  xnor keyGate_0_43(KeyNOTWire_0[24], keyinput43, keyinput_Wire_0[43]);
  not KeyNOTGate_0_24(N321, KeyNOTWire_0[24]);
  xor XOR2_57 (keyinput_Wire_0[44], N290, N293);
  xnor keyGate_0_44(KeyNOTWire_0[25], keyinput44, keyinput_Wire_0[44]);
  not KeyNOTGate_0_25(N338, KeyNOTWire_0[25]);
xor XOR2_58 (N339, N296, N299);
  xor XOR2_59 (keyinput_Wire_0[45], N290, N296);
  xnor keyGate_0_45(N340, keyinput45, keyinput_Wire_0[45]);
xor XOR2_60 (N341, N293, N299);
  xor XOR2_61 (keyinput_Wire_0[46], N302, N305);
  xnor keyGate_0_46(KeyNOTWire_0[26], keyinput46, keyinput_Wire_0[46]);
  not KeyNOTGate_0_26(N342, KeyNOTWire_0[26]);
  xor XOR2_62 (keyinput_Wire_0[47], N308, N311);
  xnor keyGate_0_47(KeyNOTWire_0[27], keyinput47, keyinput_Wire_0[47]);
  not KeyNOTGate_0_27(N343, KeyNOTWire_0[27]);
  xor XOR2_63 (keyinput_Wire_0[48], N302, N308);
  xor keyGate_0_48(N344, keyinput48, keyinput_Wire_0[48]);
xor XOR2_64 (N345, N305, N311);
xor XOR2_65 (N346, N266, N342);
  xor XOR2_66 (keyinput_Wire_0[49], N267, N343);
  xor keyGate_0_49(KeyNOTWire_0[28], keyinput49, keyinput_Wire_0[49]);
  not KeyNOTGate_0_28(N347, KeyNOTWire_0[28]);
  xor XOR2_67 (keyinput_Wire_0[50], N268, N344);
  xor keyGate_0_50(N348, keyinput50, keyinput_Wire_0[50]);
xor XOR2_68 (N349, N269, N345);
  xor XOR2_69 (keyinput_Wire_0[51], N270, N338);
  xnor keyGate_0_51(KeyNOTWire_0[29], keyinput51, keyinput_Wire_0[51]);
  not KeyNOTGate_0_29(N350, KeyNOTWire_0[29]);
  xor XOR2_70 (keyinput_Wire_0[52], N271, N339);
  xor keyGate_0_52(N351, keyinput52, keyinput_Wire_0[52]);
  xor XOR2_71 (keyinput_Wire_0[53], N272, N340);
  xor keyGate_0_53(N352, keyinput53, keyinput_Wire_0[53]);
  xor XOR2_72 (keyinput_Wire_0[54], N273, N341);
  xor keyGate_0_54(N353, keyinput54, keyinput_Wire_0[54]);
  xor XOR2_73 (keyinput_Wire_0[55], N314, N346);
  xnor keyGate_0_55(N354, keyinput55, keyinput_Wire_0[55]);
  xor XOR2_74 (keyinput_Wire_0[56], N315, N347);
  xor keyGate_0_56(KeyNOTWire_0[30], keyinput56, keyinput_Wire_0[56]);
  not KeyNOTGate_0_30(N367, KeyNOTWire_0[30]);
  xor XOR2_75 (keyinput_Wire_0[57], N316, N348);
  xor keyGate_0_57(N380, keyinput57, keyinput_Wire_0[57]);
xor XOR2_76 (N393, N317, N349);
xor XOR2_77 (N406, N318, N350);
  xor XOR2_78 (keyinput_Wire_0[58], N319, N351);
  xor keyGate_0_58(N419, keyinput58, keyinput_Wire_0[58]);
xor XOR2_79 (N432, N320, N352);
xor XOR2_80 (N445, N321, N353);
not NOT1_81 (N554, N354);
not NOT1_82 (N555, N367);
not NOT1_83 (N556, N380);
not NOT1_84 (N557, N354);
not NOT1_85 (N558, N367);
not NOT1_86 (N559, N393);
not NOT1_87 (N560, N354);
not NOT1_88 (N561, N380);
not NOT1_89 (N562, N393);
not NOT1_90 (N563, N367);
not NOT1_91 (N564, N380);
not NOT1_92 (N565, N393);
not NOT1_93 (N566, N419);
not NOT1_94 (N567, N445);
not NOT1_95 (N568, N419);
not NOT1_96 (N569, N432);
not NOT1_97 (N570, N406);
not NOT1_98 (N571, N445);
not NOT1_99 (N572, N406);
not NOT1_100 (N573, N432);
not NOT1_101 (N574, N406);
not NOT1_102 (N575, N419);
not NOT1_103 (N576, N432);
not NOT1_104 (N577, N406);
not NOT1_105 (N578, N419);
not NOT1_106 (N579, N445);
not NOT1_107 (N580, N406);
not NOT1_108 (N581, N432);
not NOT1_109 (N582, N445);
not NOT1_110 (N583, N419);
not NOT1_111 (N584, N432);
not NOT1_112 (N585, N445);
not NOT1_113 (N586, N367);
not NOT1_114 (N587, N393);
not NOT1_115 (N588, N367);
not NOT1_116 (N589, N380);
not NOT1_117 (N590, N354);
not NOT1_118 (N591, N393);
not NOT1_119 (N592, N354);
not NOT1_120 (N593, N380);
and AND4_121 (N594, N554, N555, N556, N393);
and AND4_122 (N595, N557, N558, N380, N559);
and AND4_123 (N596, N560, N367, N561, N562);
and AND4_124 (N597, N354, N563, N564, N565);
and AND4_125 (N598, N574, N575, N576, N445);
and AND4_126 (N599, N577, N578, N432, N579);
and AND4_127 (N600, N580, N419, N581, N582);
and AND4_128 (N601, N406, N583, N584, N585);
or OR4_129 (N602, N594, N595, N596, N597);
or OR4_130 (N607, N598, N599, N600, N601);
and AND5_131 (N620, N406, N566, N432, N567, N602);
and AND5_132 (N625, N406, N568, N569, N445, N602);
and AND5_133 (N630, N570, N419, N432, N571, N602);
and AND5_134 (N635, N572, N419, N573, N445, N602);
and AND5_135 (N640, N354, N586, N380, N587, N607);
  and AND5_136 (keyinput_Wire_0[59], N354, N588, N589, N393, N607);
  xnor keyGate_0_59(KeyNOTWire_0[31], keyinput59, keyinput_Wire_0[59]);
  not KeyNOTGate_0_31(N645, KeyNOTWire_0[31]);
and AND5_137 (N650, N590, N367, N380, N591, N607);
and AND5_138 (N655, N592, N367, N593, N393, N607);
and AND2_139 (N692, N354, N620);
and AND2_140 (N693, N367, N620);
and AND2_141 (N694, N380, N620);
and AND2_142 (N695, N393, N620);
and AND2_143 (N696, N354, N625);
and AND2_144 (N697, N367, N625);
and AND2_145 (N698, N380, N625);
and AND2_146 (N699, N393, N625);
and AND2_147 (N700, N354, N630);
and AND2_148 (N701, N367, N630);
and AND2_149 (N702, N380, N630);
and AND2_150 (N703, N393, N630);
and AND2_151 (N704, N354, N635);
and AND2_152 (N705, N367, N635);
and AND2_153 (N706, N380, N635);
  and AND2_154 (keyinput_Wire_0[60], N393, N635);
  xor keyGate_0_60(N707, keyinput60, keyinput_Wire_0[60]);
and AND2_155 (N708, N406, N640);
and AND2_156 (N709, N419, N640);
and AND2_157 (N710, N432, N640);
and AND2_158 (N711, N445, N640);
and AND2_159 (N712, N406, N645);
  and AND2_160 (keyinput_Wire_0[61], N419, N645);
  xor keyGate_0_61(KeyNOTWire_0[32], keyinput61, keyinput_Wire_0[61]);
  not KeyNOTGate_0_32(N713, KeyNOTWire_0[32]);
and AND2_161 (N714, N432, N645);
  and AND2_162 (keyinput_Wire_0[62], N445, N645);
  xnor keyGate_0_62(N715, keyinput62, keyinput_Wire_0[62]);
and AND2_163 (N716, N406, N650);
and AND2_164 (N717, N419, N650);
and AND2_165 (N718, N432, N650);
and AND2_166 (N719, N445, N650);
and AND2_167 (N720, N406, N655);
and AND2_168 (N721, N419, N655);
and AND2_169 (N722, N432, N655);
and AND2_170 (N723, N445, N655);
xor XOR2_171 (N724, N1, N692);
xor XOR2_172 (N725, N5, N693);
xor XOR2_173 (N726, N9, N694);
xor XOR2_174 (N727, N13, N695);
xor XOR2_175 (N728, N17, N696);
xor XOR2_176 (N729, N21, N697);
xor XOR2_177 (N730, N25, N698);
xor XOR2_178 (N731, N29, N699);
xor XOR2_179 (N732, N33, N700);
xor XOR2_180 (N733, N37, N701);
xor XOR2_181 (N734, N41, N702);
xor XOR2_182 (N735, N45, N703);
xor XOR2_183 (N736, N49, N704);
xor XOR2_184 (N737, N53, N705);
xor XOR2_185 (N738, N57, N706);
xor XOR2_186 (N739, N61, N707);
xor XOR2_187 (KeyWire_0_1, N65, N708);
  xor flip_it (N740, KeyWire_0_1, KeyWire_0_2 );
xor XOR2_188 (N741, N69, N709);
xor XOR2_189 (N742, N73, N710);
xor XOR2_190 (N743, N77, N711);
xor XOR2_191 (N744, N81, N712);
xor XOR2_192 (N745, N85, N713);
  xor XOR2_193 (keyinput_Wire_0[63], N89, N714);
  xnor keyGate_0_63(N746, keyinput63, keyinput_Wire_0[63]);
xor XOR2_194 (N747, N93, N715);
xor XOR2_195 (N748, N97, N716);
xor XOR2_196 (N749, N101, N717);
xor XOR2_197 (N750, N105, N718);
xor XOR2_198 (N751, N109, N719);
xor XOR2_199 (N752, N113, N720);
xor XOR2_200 (N753, N117, N721);
xor XOR2_201 (N754, N121, N722);
xor XOR2_202 (N755, N125, N723);

AntiSAT some_name( KeyWire_0_2, N135, N65, N13, N89, N41, N5, N93, N109, N17, N9, N136, N61, N117, N53, N33, N29, N49, N125, N113, N105, N37, N101, N130, N134, N137, N133, N81, N85, N129, N97, N132, N45, N1, N21, N69, N131, N57, N73, N77, N121, N25, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145,
       keyinput146, keyinput147, keyinput148, keyinput149, keyinput150,
       keyinput151, keyinput152, keyinput153, keyinput154, keyinput155,
       keyinput156, keyinput157, keyinput158, keyinput159, keyinput160,
       keyinput161, keyinput162, keyinput163, keyinput164, keyinput165,
       keyinput166, keyinput167, keyinput168, keyinput169, keyinput170,
       keyinput171, keyinput172, keyinput173, keyinput174, keyinput175,
       keyinput176, keyinput177, keyinput178, keyinput179, keyinput180,
       keyinput181, keyinput182, keyinput183, keyinput184, keyinput185,
       keyinput186);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N135, N65, N13, N89, N41, N5, N93, N109, N17, N9, N136, N61, N117, N53, N33, N29, N49, N125, N113, N105, N37, N101, N130, N134, N137, N133, N81, N85, N129, N97, N132, N45, N1, N21, N69, N131, N57, N73, N77, N121, N25, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145 ,
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150,
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155,
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160,
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165,
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170,
        keyinput171, keyinput172, keyinput173, keyinput174, keyinput175,
        keyinput176, keyinput177, keyinput178, keyinput179, keyinput180,
        keyinput181, keyinput182, keyinput183, keyinput184, keyinput185,
        keyinput186);

  input keyinput146, keyinput147, keyinput148, keyinput149, keyinput150;
  input keyinput151, keyinput152, keyinput153, keyinput154, keyinput155;
  input keyinput156, keyinput157, keyinput158, keyinput159, keyinput160;
  input keyinput161, keyinput162, keyinput163, keyinput164, keyinput165;
  input keyinput166, keyinput167, keyinput168, keyinput169, keyinput170;
  input keyinput171, keyinput172, keyinput173, keyinput174, keyinput175;
  input keyinput176, keyinput177, keyinput178, keyinput179, keyinput180;
  input keyinput181, keyinput182, keyinput183, keyinput184, keyinput185;
  input keyinput186;

  wire [0:40] keyNTin_Wire_1;
  wire [0:19] KeyNOTWire_1;

  input N135, N65, N13, N89, N41, N5, N93, N109, N17, N9, N136, N61, N117, N53, N33, N29, N49, N125, N113, N105, N37, N101, N130, N134, N137, N133, N81, N85, N129, N97, N132, N45, N1, N21, N69, N131, N57, N73, N77, N121, N25;
  input keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, keyinput145;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83 ;

  xnor KeyGate0 (newWire_0, N135, keyinput64);
  xnor KeyGate1 (newWire_1, N65, keyinput65);
  xnor KeyGate2 (newWire_2, N13, keyinput66);
  xor  KeyGate3 (keyNTin_Wire_1[0], N89, keyinput67);
  xnor keyNTinGate_1_0(KeyNOTWire_1[0], keyinput146, keyNTin_Wire_1[0]);
  not KeyNOTGate_1_0(newWire_3, KeyNOTWire_1[0]);
  xnor KeyGate4 (newWire_4, N41, keyinput68);
  xnor KeyGate5 (keyNTin_Wire_1[1], N5, keyinput69);
  xnor keyNTinGate_1_1(KeyNOTWire_1[1], keyinput147, keyNTin_Wire_1[1]);
  not KeyNOTGate_1_1(newWire_5, KeyNOTWire_1[1]);
  xor  KeyGate6 (keyNTin_Wire_1[2], N93, keyinput70);
  xor keyNTinGate_1_2(KeyNOTWire_1[2], keyinput148, keyNTin_Wire_1[2]);
  not KeyNOTGate_1_2(newWire_6, KeyNOTWire_1[2]);
  xnor KeyGate7 (keyNTin_Wire_1[3], N109, keyinput71);
  xnor keyNTinGate_1_3(newWire_7, keyinput149, keyNTin_Wire_1[3]);
  xor  KeyGate8 (newWire_8, N17, keyinput72);
  xor  KeyGate9 (newWire_9, N9, keyinput73);
  xor  KeyGate10 (newWire_10, N136, keyinput74);
  xnor KeyGate11 (newWire_11, N61, keyinput75);
  xor  KeyGate12 (newWire_12, N117, keyinput76);
  xor  KeyGate13 (newWire_13, N53, keyinput77);
  xnor KeyGate14 (keyNTin_Wire_1[4], N33, keyinput78);
  xor keyNTinGate_1_4(KeyNOTWire_1[3], keyinput150, keyNTin_Wire_1[4]);
  not KeyNOTGate_1_3(newWire_14, KeyNOTWire_1[3]);
  xor  KeyGate15 (keyNTin_Wire_1[5], N29, keyinput79);
  xor keyNTinGate_1_5(newWire_15, keyinput151, keyNTin_Wire_1[5]);
  xnor KeyGate16 (newWire_16, N49, keyinput80);
  xor  KeyGate17 (keyNTin_Wire_1[6], N125, keyinput81);
  xor keyNTinGate_1_6(KeyNOTWire_1[4], keyinput152, keyNTin_Wire_1[6]);
  not KeyNOTGate_1_4(newWire_17, KeyNOTWire_1[4]);
  xnor KeyGate18 (newWire_18, N113, keyinput82);
  xor  KeyGate19 (newWire_19, N105, keyinput83);
  xor  KeyGate20 (keyNTin_Wire_1[7], N37, keyinput84);
  xor keyNTinGate_1_7(KeyNOTWire_1[5], keyinput153, keyNTin_Wire_1[7]);
  not KeyNOTGate_1_5(newWire_20, KeyNOTWire_1[5]);
  xnor KeyGate21 (keyNTin_Wire_1[8], N101, keyinput85);
  xnor keyNTinGate_1_8(KeyNOTWire_1[6], keyinput154, keyNTin_Wire_1[8]);
  not KeyNOTGate_1_6(newWire_21, KeyNOTWire_1[6]);
  xnor KeyGate22 (keyNTin_Wire_1[9], N130, keyinput86);
  xnor keyNTinGate_1_9(KeyNOTWire_1[7], keyinput155, keyNTin_Wire_1[9]);
  not KeyNOTGate_1_7(newWire_22, KeyNOTWire_1[7]);
  xor  KeyGate23 (newWire_23, N134, keyinput87);
  xnor KeyGate24 (newWire_24, N137, keyinput88);
  xnor KeyGate25 (keyNTin_Wire_1[10], N133, keyinput89);
  xnor keyNTinGate_1_10(KeyNOTWire_1[8], keyinput156, keyNTin_Wire_1[10]);
  not KeyNOTGate_1_8(newWire_25, KeyNOTWire_1[8]);
  xnor KeyGate26 (newWire_26, N81, keyinput90);
  xor  KeyGate27 (keyNTin_Wire_1[11], N85, keyinput91);
  xnor keyNTinGate_1_11(KeyNOTWire_1[9], keyinput157, keyNTin_Wire_1[11]);
  not KeyNOTGate_1_9(newWire_27, KeyNOTWire_1[9]);
  xnor KeyGate28 (keyNTin_Wire_1[12], N129, keyinput92);
  xor keyNTinGate_1_12(newWire_28, keyinput158, keyNTin_Wire_1[12]);
  xor  KeyGate29 (keyNTin_Wire_1[13], N97, keyinput93);
  xnor keyNTinGate_1_13(newWire_29, keyinput159, keyNTin_Wire_1[13]);
  xor  KeyGate30 (newWire_30, N132, keyinput94);
  xor  KeyGate31 (keyNTin_Wire_1[14], N45, keyinput95);
  xnor keyNTinGate_1_14(KeyNOTWire_1[10], keyinput160, keyNTin_Wire_1[14]);
  not KeyNOTGate_1_10(newWire_31, KeyNOTWire_1[10]);
  xnor KeyGate32 (keyNTin_Wire_1[15], N1, keyinput96);
  xor keyNTinGate_1_15(newWire_32, keyinput161, keyNTin_Wire_1[15]);
  xnor KeyGate33 (newWire_33, N21, keyinput97);
  xnor KeyGate34 (newWire_34, N69, keyinput98);
  xor  KeyGate35 (keyNTin_Wire_1[16], N131, keyinput99);
  xor keyNTinGate_1_16(KeyNOTWire_1[11], keyinput162, keyNTin_Wire_1[16]);
  not KeyNOTGate_1_11(newWire_35, KeyNOTWire_1[11]);
  xor  KeyGate36 (keyNTin_Wire_1[17], N57, keyinput100);
  xor keyNTinGate_1_17(newWire_36, keyinput163, keyNTin_Wire_1[17]);
  xnor KeyGate37 (newWire_37, N73, keyinput101);
  xor  KeyGate38 (newWire_38, N77, keyinput102);
  xnor KeyGate39 (newWire_39, N121, keyinput103);
  xnor KeyGate40 (newWire_40, N25, keyinput104);
  xnor KeyGate41 (keyNTin_Wire_1[18], N135, keyinput105);
  xor keyNTinGate_1_18(newWire_41, keyinput164, keyNTin_Wire_1[18]);
  xor  KeyGate42 (newWire_42, N65, keyinput106);
  xnor KeyGate43 (keyNTin_Wire_1[19], N13, keyinput107);
  xor keyNTinGate_1_19(KeyNOTWire_1[12], keyinput165, keyNTin_Wire_1[19]);
  not KeyNOTGate_1_12(newWire_43, KeyNOTWire_1[12]);
  xnor KeyGate44 (newWire_44, N89, keyinput108);
  xnor KeyGate45 (keyNTin_Wire_1[20], N41, keyinput109);
  xnor keyNTinGate_1_20(newWire_45, keyinput166, keyNTin_Wire_1[20]);
  xnor KeyGate46 (newWire_46, N5, keyinput110);
  xor  KeyGate47 (newWire_47, N93, keyinput111);
  xnor KeyGate48 (newWire_48, N109, keyinput112);
  xnor KeyGate49 (newWire_49, N17, keyinput113);
  xor  KeyGate50 (keyNTin_Wire_1[21], N9, keyinput114);
  xnor keyNTinGate_1_21(newWire_50, keyinput167, keyNTin_Wire_1[21]);
  xor  KeyGate51 (newWire_51, N136, keyinput115);
  xnor KeyGate52 (keyNTin_Wire_1[22], N61, keyinput116);
  xnor keyNTinGate_1_22(newWire_52, keyinput168, keyNTin_Wire_1[22]);
  xor  KeyGate53 (newWire_53, N117, keyinput117);
  xnor KeyGate54 (keyNTin_Wire_1[23], N53, keyinput118);
  xor keyNTinGate_1_23(KeyNOTWire_1[13], keyinput169, keyNTin_Wire_1[23]);
  not KeyNOTGate_1_13(newWire_54, KeyNOTWire_1[13]);
  xor  KeyGate55 (newWire_55, N33, keyinput119);
  xnor KeyGate56 (keyNTin_Wire_1[24], N29, keyinput120);
  xor keyNTinGate_1_24(KeyNOTWire_1[14], keyinput170, keyNTin_Wire_1[24]);
  not KeyNOTGate_1_14(newWire_56, KeyNOTWire_1[14]);
  xnor KeyGate57 (newWire_57, N49, keyinput121);
  xnor KeyGate58 (keyNTin_Wire_1[25], N125, keyinput122);
  xor keyNTinGate_1_25(newWire_58, keyinput171, keyNTin_Wire_1[25]);
  xnor KeyGate59 (newWire_59, N113, keyinput123);
  xor  KeyGate60 (keyNTin_Wire_1[26], N105, keyinput124);
  xor keyNTinGate_1_26(newWire_60, keyinput172, keyNTin_Wire_1[26]);
  xnor KeyGate61 (keyNTin_Wire_1[27], N37, keyinput125);
  xor keyNTinGate_1_27(KeyNOTWire_1[15], keyinput173, keyNTin_Wire_1[27]);
  not KeyNOTGate_1_15(newWire_61, KeyNOTWire_1[15]);
  xor  KeyGate62 (keyNTin_Wire_1[28], N101, keyinput126);
  xor keyNTinGate_1_28(newWire_62, keyinput174, keyNTin_Wire_1[28]);
  xnor KeyGate63 (newWire_63, N130, keyinput127);
  xnor KeyGate64 (keyNTin_Wire_1[29], N134, keyinput128);
  xnor keyNTinGate_1_29(newWire_64, keyinput175, keyNTin_Wire_1[29]);
  xnor KeyGate65 (keyNTin_Wire_1[30], N137, keyinput129);
  xnor keyNTinGate_1_30(KeyNOTWire_1[16], keyinput176, keyNTin_Wire_1[30]);
  not KeyNOTGate_1_16(newWire_65, KeyNOTWire_1[16]);
  xnor KeyGate66 (newWire_66, N133, keyinput130);
  xnor KeyGate67 (newWire_67, N81, keyinput131);
  xnor KeyGate68 (keyNTin_Wire_1[31], N85, keyinput132);
  xor keyNTinGate_1_31(newWire_68, keyinput177, keyNTin_Wire_1[31]);
  xnor KeyGate69 (keyNTin_Wire_1[32], N129, keyinput133);
  xor keyNTinGate_1_32(KeyNOTWire_1[17], keyinput178, keyNTin_Wire_1[32]);
  not KeyNOTGate_1_17(newWire_69, KeyNOTWire_1[17]);
  xnor KeyGate70 (newWire_70, N97, keyinput134);
  xnor KeyGate71 (keyNTin_Wire_1[33], N132, keyinput135);
  xor keyNTinGate_1_33(newWire_71, keyinput179, keyNTin_Wire_1[33]);
  xor  KeyGate72 (keyNTin_Wire_1[34], N45, keyinput136);
  xor keyNTinGate_1_34(KeyNOTWire_1[18], keyinput180, keyNTin_Wire_1[34]);
  not KeyNOTGate_1_18(newWire_72, KeyNOTWire_1[18]);
  xnor KeyGate73 (keyNTin_Wire_1[35], N1, keyinput137);
  xnor keyNTinGate_1_35(newWire_73, keyinput181, keyNTin_Wire_1[35]);
  xor  KeyGate74 (keyNTin_Wire_1[36], N21, keyinput138);
  xor keyNTinGate_1_36(newWire_74, keyinput182, keyNTin_Wire_1[36]);
  xnor KeyGate75 (newWire_75, N69, keyinput139);
  xor  KeyGate76 (keyNTin_Wire_1[37], N131, keyinput140);
  xor keyNTinGate_1_37(newWire_76, keyinput183, keyNTin_Wire_1[37]);
  xor  KeyGate77 (keyNTin_Wire_1[38], N57, keyinput141);
  xnor keyNTinGate_1_38(KeyNOTWire_1[19], keyinput184, keyNTin_Wire_1[38]);
  not KeyNOTGate_1_19(newWire_77, KeyNOTWire_1[19]);
  xnor KeyGate78 (newWire_78, N73, keyinput142);
  xor  KeyGate79 (newWire_79, N77, keyinput143);
  xnor KeyGate80 (keyNTin_Wire_1[39], N121, keyinput144);
  xnor keyNTinGate_1_39(newWire_80, keyinput185, keyNTin_Wire_1[39]);
  xnor KeyGate81 (newWire_81, N25, keyinput145);
  and some_function (newWire_82, newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40 );
  nand compl_function (keyNTin_Wire_1[40], newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81);
  xor keyNTinGate_1_40(newWire_83, keyinput186, keyNTin_Wire_1[40]);
  and finalAND (KeyWire_0_2, newWire_82, newWire_83);

endmodule /* AntiSAT */
