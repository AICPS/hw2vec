`timescale 1ns / 1ps
// Verilog
// c499
// Ninputs 41
// Noutputs 32
// NtotalGates 202
// XOR2 104
// AND2 40
// NOT1 40
// AND4 8
// OR4 2
// AND5 8

module top (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
                  N753,N754,N755,
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
                  keyinput30, keyinput31,
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36,
        keyinput37, keyinput38, keyinput39, keyinput40, keyinput41,
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46,
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51,
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56,
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61,
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66,
        keyinput67, keyinput68, keyinput69, keyinput70, keyinput71,
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76,
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81,
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86,
        keyinput87, keyinput88, keyinput89, keyinput90, keyinput91,
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96,
        keyinput97, keyinput98, keyinput99, keyinput100, keyinput101,
        keyinput102, keyinput103, keyinput104, keyinput105, keyinput106,
        keyinput107, keyinput108, keyinput109, keyinput110, keyinput111,
                  keyinput112, keyinput113,
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
        keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
        keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
        keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
        keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
        keyinput144, keyinput145, keyinput146, keyinput147, keyinput148,
        keyinput149, keyinput150, keyinput151, keyinput152, keyinput153,
        keyinput154);

  input keyinput114, keyinput115, keyinput116, keyinput117, keyinput118;
  input keyinput119, keyinput120, keyinput121, keyinput122, keyinput123;
  input keyinput124, keyinput125, keyinput126, keyinput127, keyinput128;
  input keyinput129, keyinput130, keyinput131, keyinput132, keyinput133;
  input keyinput134, keyinput135, keyinput136, keyinput137, keyinput138;
  input keyinput139, keyinput140, keyinput141, keyinput142, keyinput143;
  input keyinput144, keyinput145, keyinput146, keyinput147, keyinput148;
  input keyinput149, keyinput150, keyinput151, keyinput152, keyinput153;
  input keyinput154;


  input keyinput32, keyinput33, keyinput34, keyinput35, keyinput36;
  input keyinput37, keyinput38, keyinput39, keyinput40, keyinput41;
  input keyinput42, keyinput43, keyinput44, keyinput45, keyinput46;
  input keyinput47, keyinput48, keyinput49, keyinput50, keyinput51;
  input keyinput52, keyinput53, keyinput54, keyinput55, keyinput56;
  input keyinput57, keyinput58, keyinput59, keyinput60, keyinput61;
  input keyinput62, keyinput63, keyinput64, keyinput65, keyinput66;
  input keyinput67, keyinput68, keyinput69, keyinput70, keyinput71;
  input keyinput72, keyinput73, keyinput74, keyinput75, keyinput76;
  input keyinput77, keyinput78, keyinput79, keyinput80, keyinput81;
  input keyinput82, keyinput83, keyinput84, keyinput85, keyinput86;
  input keyinput87, keyinput88, keyinput89, keyinput90, keyinput91;
  input keyinput92, keyinput93, keyinput94, keyinput95, keyinput96;
  input keyinput97, keyinput98, keyinput99, keyinput100, keyinput101;
  input keyinput102, keyinput103, keyinput104, keyinput105, keyinput106;
  input keyinput107, keyinput108, keyinput109, keyinput110, keyinput111;
  input keyinput112, keyinput113;

  wire KeyWire_0_1 , KeyWire_0_2;

  input keyinput0, keyinput1, keyinput2, keyinput3, keyinput4;
  input keyinput5, keyinput6, keyinput7, keyinput8, keyinput9;
  input keyinput10, keyinput11, keyinput12, keyinput13, keyinput14;
  input keyinput15, keyinput16, keyinput17, keyinput18, keyinput19;
  input keyinput20, keyinput21, keyinput22, keyinput23, keyinput24;
  input keyinput25, keyinput26, keyinput27, keyinput28, keyinput29;
  input keyinput30, keyinput31;

  wire [0:31] keyinput_Wire_0;
  wire [0:13] KeyNOTWire_0;

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;

output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723;

  xor XOR2_1 (keyinput_Wire_0[0], N1, N5);
  xor keyGate_0_0(N250, keyinput0, keyinput_Wire_0[0]);
  xor XOR2_2 (keyinput_Wire_0[1], N9, N13);
  xor keyGate_0_1(N251, keyinput1, keyinput_Wire_0[1]);
  xor XOR2_3 (keyinput_Wire_0[2], N17, N21);
  xnor keyGate_0_2(KeyNOTWire_0[0], keyinput2, keyinput_Wire_0[2]);
  not KeyNOTGate_0_0(N252, KeyNOTWire_0[0]);
  xor XOR2_4 (keyinput_Wire_0[3], N25, N29);
  xnor keyGate_0_3(KeyNOTWire_0[1], keyinput3, keyinput_Wire_0[3]);
  not KeyNOTGate_0_1(N253, KeyNOTWire_0[1]);
  xor XOR2_5 (keyinput_Wire_0[4], N33, N37);
  xnor keyGate_0_4(N254, keyinput4, keyinput_Wire_0[4]);
  xor XOR2_6 (keyinput_Wire_0[5], N41, N45);
  xor keyGate_0_5(N255, keyinput5, keyinput_Wire_0[5]);
  xor XOR2_7 (keyinput_Wire_0[6], N49, N53);
  xor keyGate_0_6(KeyNOTWire_0[2], keyinput6, keyinput_Wire_0[6]);
  not KeyNOTGate_0_2(N256, KeyNOTWire_0[2]);
  xor XOR2_8 (keyinput_Wire_0[7], N57, N61);
  xnor keyGate_0_7(N257, keyinput7, keyinput_Wire_0[7]);
  xor XOR2_9 (keyinput_Wire_0[8], N65, N69);
  xor keyGate_0_8(N258, keyinput8, keyinput_Wire_0[8]);
xor XOR2_10 (N259, N73, N77);
xor XOR2_11 (N260, N81, N85);
xor XOR2_12 (N261, N89, N93);
xor XOR2_13 (N262, N97, N101);
xor XOR2_14 (N263, N105, N109);
xor XOR2_15 (N264, N113, N117);
xor XOR2_16 (N265, N121, N125);
and AND2_17 (N266, N129, N137);
and AND2_18 (N267, N130, N137);
and AND2_19 (N268, N131, N137);
and AND2_20 (N269, N132, N137);
and AND2_21 (N270, N133, N137);
and AND2_22 (N271, N134, N137);
and AND2_23 (N272, N135, N137);
and AND2_24 (N273, N136, N137);
xor XOR2_25 (N274, N1, N17);
xor XOR2_26 (N275, N33, N49);
xor XOR2_27 (N276, N5, N21);
xor XOR2_28 (N277, N37, N53);
xor XOR2_29 (N278, N9, N25);
xor XOR2_30 (N279, N41, N57);
xor XOR2_31 (N280, N13, N29);
xor XOR2_32 (N281, N45, N61);
xor XOR2_33 (N282, N65, N81);
xor XOR2_34 (N283, N97, N113);
xor XOR2_35 (N284, N69, N85);
xor XOR2_36 (N285, N101, N117);
xor XOR2_37 (N286, N73, N89);
xor XOR2_38 (N287, N105, N121);
xor XOR2_39 (N288, N77, N93);
xor XOR2_40 (N289, N109, N125);
  xor XOR2_41 (keyinput_Wire_0[9], N250, N251);
  xor keyGate_0_9(N290, keyinput9, keyinput_Wire_0[9]);
  xor XOR2_42 (keyinput_Wire_0[10], N252, N253);
  xor keyGate_0_10(KeyNOTWire_0[3], keyinput10, keyinput_Wire_0[10]);
  not KeyNOTGate_0_3(N293, KeyNOTWire_0[3]);
  xor XOR2_43 (keyinput_Wire_0[11], N254, N255);
  xor keyGate_0_11(N296, keyinput11, keyinput_Wire_0[11]);
  xor XOR2_44 (keyinput_Wire_0[12], N256, N257);
  xor keyGate_0_12(KeyNOTWire_0[4], keyinput12, keyinput_Wire_0[12]);
  not KeyNOTGate_0_4(N299, KeyNOTWire_0[4]);
  xor XOR2_45 (keyinput_Wire_0[13], N258, N259);
  xor keyGate_0_13(N302, keyinput13, keyinput_Wire_0[13]);
  xor XOR2_46 (keyinput_Wire_0[14], N260, N261);
  xnor keyGate_0_14(KeyNOTWire_0[5], keyinput14, keyinput_Wire_0[14]);
  not KeyNOTGate_0_5(N305, KeyNOTWire_0[5]);
  xor XOR2_47 (keyinput_Wire_0[15], N262, N263);
  xor keyGate_0_15(KeyNOTWire_0[6], keyinput15, keyinput_Wire_0[15]);
  not KeyNOTGate_0_6(N308, KeyNOTWire_0[6]);
  xor XOR2_48 (keyinput_Wire_0[16], N264, N265);
  xor keyGate_0_16(N311, keyinput16, keyinput_Wire_0[16]);
xor XOR2_49 (N314, N274, N275);
xor XOR2_50 (N315, N276, N277);
xor XOR2_51 (N316, N278, N279);
xor XOR2_52 (N317, N280, N281);
xor XOR2_53 (N318, N282, N283);
xor XOR2_54 (N319, N284, N285);
xor XOR2_55 (N320, N286, N287);
xor XOR2_56 (N321, N288, N289);
xor XOR2_57 (N338, N290, N293);
xor XOR2_58 (N339, N296, N299);
xor XOR2_59 (N340, N290, N296);
xor XOR2_60 (N341, N293, N299);
xor XOR2_61 (N342, N302, N305);
xor XOR2_62 (N343, N308, N311);
xor XOR2_63 (N344, N302, N308);
xor XOR2_64 (N345, N305, N311);
xor XOR2_65 (N346, N266, N342);
xor XOR2_66 (N347, N267, N343);
xor XOR2_67 (N348, N268, N344);
xor XOR2_68 (N349, N269, N345);
xor XOR2_69 (N350, N270, N338);
xor XOR2_70 (N351, N271, N339);
xor XOR2_71 (N352, N272, N340);
xor XOR2_72 (N353, N273, N341);
xor XOR2_73 (N354, N314, N346);
xor XOR2_74 (N367, N315, N347);
xor XOR2_75 (N380, N316, N348);
xor XOR2_76 (N393, N317, N349);
xor XOR2_77 (N406, N318, N350);
xor XOR2_78 (N419, N319, N351);
xor XOR2_79 (N432, N320, N352);
xor XOR2_80 (N445, N321, N353);
not NOT1_81 (N554, N354);
not NOT1_82 (N555, N367);
not NOT1_83 (N556, N380);
not NOT1_84 (N557, N354);
not NOT1_85 (N558, N367);
not NOT1_86 (N559, N393);
not NOT1_87 (N560, N354);
not NOT1_88 (N561, N380);
not NOT1_89 (N562, N393);
not NOT1_90 (N563, N367);
not NOT1_91 (N564, N380);
not NOT1_92 (N565, N393);
not NOT1_93 (N566, N419);
not NOT1_94 (N567, N445);
not NOT1_95 (N568, N419);
not NOT1_96 (N569, N432);
not NOT1_97 (N570, N406);
not NOT1_98 (N571, N445);
not NOT1_99 (N572, N406);
not NOT1_100 (N573, N432);
not NOT1_101 (N574, N406);
not NOT1_102 (N575, N419);
not NOT1_103 (N576, N432);
not NOT1_104 (N577, N406);
not NOT1_105 (N578, N419);
not NOT1_106 (N579, N445);
not NOT1_107 (N580, N406);
not NOT1_108 (N581, N432);
not NOT1_109 (N582, N445);
not NOT1_110 (N583, N419);
not NOT1_111 (N584, N432);
not NOT1_112 (N585, N445);
not NOT1_113 (N586, N367);
not NOT1_114 (N587, N393);
not NOT1_115 (N588, N367);
not NOT1_116 (N589, N380);
not NOT1_117 (N590, N354);
not NOT1_118 (N591, N393);
not NOT1_119 (N592, N354);
not NOT1_120 (N593, N380);
and AND4_121 (N594, N554, N555, N556, N393);
and AND4_122 (N595, N557, N558, N380, N559);
and AND4_123 (N596, N560, N367, N561, N562);
and AND4_124 (N597, N354, N563, N564, N565);
and AND4_125 (N598, N574, N575, N576, N445);
and AND4_126 (N599, N577, N578, N432, N579);
and AND4_127 (N600, N580, N419, N581, N582);
and AND4_128 (N601, N406, N583, N584, N585);
or OR4_129 (N602, N594, N595, N596, N597);
or OR4_130 (N607, N598, N599, N600, N601);
  and AND5_131 (keyinput_Wire_0[17], N406, N566, N432, N567, N602);
  xnor keyGate_0_17(KeyNOTWire_0[7], keyinput17, keyinput_Wire_0[17]);
  not KeyNOTGate_0_7(N620, KeyNOTWire_0[7]);
  and AND5_132 (keyinput_Wire_0[18], N406, N568, N569, N445, N602);
  xnor keyGate_0_18(KeyNOTWire_0[8], keyinput18, keyinput_Wire_0[18]);
  not KeyNOTGate_0_8(N625, KeyNOTWire_0[8]);
  and AND5_133 (keyinput_Wire_0[19], N570, N419, N432, N571, N602);
  xnor keyGate_0_19(N630, keyinput19, keyinput_Wire_0[19]);
  and AND5_134 (keyinput_Wire_0[20], N572, N419, N573, N445, N602);
  xor keyGate_0_20(N635, keyinput20, keyinput_Wire_0[20]);
  and AND5_135 (keyinput_Wire_0[21], N354, N586, N380, N587, N607);
  xor keyGate_0_21(N640, keyinput21, keyinput_Wire_0[21]);
  and AND5_136 (keyinput_Wire_0[22], N354, N588, N589, N393, N607);
  xnor keyGate_0_22(N645, keyinput22, keyinput_Wire_0[22]);
  and AND5_137 (keyinput_Wire_0[23], N590, N367, N380, N591, N607);
  xor keyGate_0_23(N650, keyinput23, keyinput_Wire_0[23]);
  and AND5_138 (keyinput_Wire_0[24], N592, N367, N593, N393, N607);
  xnor keyGate_0_24(KeyNOTWire_0[9], keyinput24, keyinput_Wire_0[24]);
  not KeyNOTGate_0_9(N655, KeyNOTWire_0[9]);
and AND2_139 (N692, N354, N620);
and AND2_140 (N693, N367, N620);
and AND2_141 (N694, N380, N620);
and AND2_142 (N695, N393, N620);
and AND2_143 (N696, N354, N625);
and AND2_144 (N697, N367, N625);
and AND2_145 (N698, N380, N625);
and AND2_146 (N699, N393, N625);
and AND2_147 (N700, N354, N630);
and AND2_148 (N701, N367, N630);
and AND2_149 (N702, N380, N630);
and AND2_150 (N703, N393, N630);
and AND2_151 (N704, N354, N635);
and AND2_152 (N705, N367, N635);
and AND2_153 (N706, N380, N635);
and AND2_154 (N707, N393, N635);
and AND2_155 (N708, N406, N640);
and AND2_156 (N709, N419, N640);
and AND2_157 (N710, N432, N640);
and AND2_158 (N711, N445, N640);
and AND2_159 (N712, N406, N645);
and AND2_160 (N713, N419, N645);
and AND2_161 (N714, N432, N645);
and AND2_162 (N715, N445, N645);
and AND2_163 (N716, N406, N650);
and AND2_164 (N717, N419, N650);
and AND2_165 (N718, N432, N650);
and AND2_166 (N719, N445, N650);
and AND2_167 (N720, N406, N655);
and AND2_168 (N721, N419, N655);
and AND2_169 (N722, N432, N655);
and AND2_170 (N723, N445, N655);
xor XOR2_171 (N724, N1, N692);
xor XOR2_172 (N725, N5, N693);
xor XOR2_173 (N726, N9, N694);
xor XOR2_174 (N727, N13, N695);
xor XOR2_175 (N728, N17, N696);
xor XOR2_176 (N729, N21, N697);
xor XOR2_177 (N730, N25, N698);
xor XOR2_178 (N731, N29, N699);
xor XOR2_179 (N732, N33, N700);
xor XOR2_180 (N733, N37, N701);
xor XOR2_181 (N734, N41, N702);
xor XOR2_182 (N735, N45, N703);
xor XOR2_183 (N736, N49, N704);
xor XOR2_184 (N737, N53, N705);
xor XOR2_185 (N738, N57, N706);
xor XOR2_186 (N739, N61, N707);
xor XOR2_187 (N740, N65, N708);
xor XOR2_188 (N741, N69, N709);
xor XOR2_189 (N742, N73, N710);
  xor XOR2_190 (keyinput_Wire_0[25], N77, N711);
  xnor keyGate_0_25(N743, keyinput25, keyinput_Wire_0[25]);
  xor XOR2_191 (keyinput_Wire_0[26], N81, N712);
  xnor keyGate_0_26(KeyNOTWire_0[10], keyinput26, keyinput_Wire_0[26]);
  not KeyNOTGate_0_10(KeyWire_0_1, KeyNOTWire_0[10]);
  xor flip_it (N744, KeyWire_0_1, KeyWire_0_2 );
  xor XOR2_192 (keyinput_Wire_0[27], N85, N713);
  xor keyGate_0_27(KeyNOTWire_0[11], keyinput27, keyinput_Wire_0[27]);
  not KeyNOTGate_0_11(N745, KeyNOTWire_0[11]);
  xor XOR2_193 (keyinput_Wire_0[28], N89, N714);
  xor keyGate_0_28(KeyNOTWire_0[12], keyinput28, keyinput_Wire_0[28]);
  not KeyNOTGate_0_12(N746, KeyNOTWire_0[12]);
xor XOR2_194 (N747, N93, N715);
xor XOR2_195 (N748, N97, N716);
xor XOR2_196 (N749, N101, N717);
xor XOR2_197 (N750, N105, N718);
xor XOR2_198 (N751, N109, N719);
xor XOR2_199 (N752, N113, N720);
  xor XOR2_200 (keyinput_Wire_0[29], N117, N721);
  xor keyGate_0_29(KeyNOTWire_0[13], keyinput29, keyinput_Wire_0[29]);
  not KeyNOTGate_0_13(N753, KeyNOTWire_0[13]);
  xor XOR2_201 (keyinput_Wire_0[30], N121, N722);
  xnor keyGate_0_30(N754, keyinput30, keyinput_Wire_0[30]);
  xor XOR2_202 (keyinput_Wire_0[31], N125, N723);
  xnor keyGate_0_31(N755, keyinput31, keyinput_Wire_0[31]);

AntiSAT some_name( KeyWire_0_2, N49, N77, N17, N134, N129, N130, N29, N93, N65, N89, N132, N137, N136, N105, N97, N81, N101, N5, N37, N73, N1, N13, N121, N53, N69, N113, N33, N61, N9, N41, N25, N125, N131, N135, N117, N85, N57, N109, N133, N21, N45, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
       keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
       keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
       keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
       keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
       keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
       keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
       keyinput144, keyinput145, keyinput146, keyinput147, keyinput148,
       keyinput149, keyinput150, keyinput151, keyinput152, keyinput153,
       keyinput154);

endmodule

/*************************************************************************/

module AntiSAT (KeyWire_0_2, N49, N77, N17, N134, N129, N130, N29, N93, N65, N89, N132, N137, N136, N105, N97, N81, N101, N5, N37, N73, N1, N13, N121, N53, N69, N113, N33, N61, N9, N41, N25, N125, N131, N135, N117, N85, N57, N109, N133, N21, N45, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113 ,
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
        keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
        keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
        keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
        keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
        keyinput144, keyinput145, keyinput146, keyinput147, keyinput148,
        keyinput149, keyinput150, keyinput151, keyinput152, keyinput153,
        keyinput154);

  input keyinput114, keyinput115, keyinput116, keyinput117, keyinput118;
  input keyinput119, keyinput120, keyinput121, keyinput122, keyinput123;
  input keyinput124, keyinput125, keyinput126, keyinput127, keyinput128;
  input keyinput129, keyinput130, keyinput131, keyinput132, keyinput133;
  input keyinput134, keyinput135, keyinput136, keyinput137, keyinput138;
  input keyinput139, keyinput140, keyinput141, keyinput142, keyinput143;
  input keyinput144, keyinput145, keyinput146, keyinput147, keyinput148;
  input keyinput149, keyinput150, keyinput151, keyinput152, keyinput153;
  input keyinput154;

  wire [0:40] keyNTin_Wire_1;
  wire [0:21] KeyNOTWire_1;

  input N49, N77, N17, N134, N129, N130, N29, N93, N65, N89, N132, N137, N136, N105, N97, N81, N101, N5, N37, N73, N1, N13, N121, N53, N69, N113, N33, N61, N9, N41, N25, N125, N131, N135, N117, N85, N57, N109, N133, N21, N45;
  input keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, keyinput113;
  output KeyWire_0_2;
  wire newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81, newWire_82, newWire_83 ;

  xor  KeyGate0 (keyNTin_Wire_1[0], N49, keyinput32);
  xor keyNTinGate_1_0(KeyNOTWire_1[0], keyinput114, keyNTin_Wire_1[0]);
  not KeyNOTGate_1_0(newWire_0, KeyNOTWire_1[0]);
  xnor KeyGate1 (keyNTin_Wire_1[1], N77, keyinput33);
  xnor keyNTinGate_1_1(KeyNOTWire_1[1], keyinput115, keyNTin_Wire_1[1]);
  not KeyNOTGate_1_1(newWire_1, KeyNOTWire_1[1]);
  xnor KeyGate2 (keyNTin_Wire_1[2], N17, keyinput34);
  xnor keyNTinGate_1_2(newWire_2, keyinput116, keyNTin_Wire_1[2]);
  xnor KeyGate3 (keyNTin_Wire_1[3], N134, keyinput35);
  xor keyNTinGate_1_3(KeyNOTWire_1[2], keyinput117, keyNTin_Wire_1[3]);
  not KeyNOTGate_1_2(newWire_3, KeyNOTWire_1[2]);
  xor  KeyGate4 (keyNTin_Wire_1[4], N129, keyinput36);
  xnor keyNTinGate_1_4(KeyNOTWire_1[3], keyinput118, keyNTin_Wire_1[4]);
  not KeyNOTGate_1_3(newWire_4, KeyNOTWire_1[3]);
  xor  KeyGate5 (keyNTin_Wire_1[5], N130, keyinput37);
  xor keyNTinGate_1_5(KeyNOTWire_1[4], keyinput119, keyNTin_Wire_1[5]);
  not KeyNOTGate_1_4(newWire_5, KeyNOTWire_1[4]);
  xor  KeyGate6 (keyNTin_Wire_1[6], N29, keyinput38);
  xor keyNTinGate_1_6(KeyNOTWire_1[5], keyinput120, keyNTin_Wire_1[6]);
  not KeyNOTGate_1_5(newWire_6, KeyNOTWire_1[5]);
  xnor KeyGate7 (keyNTin_Wire_1[7], N93, keyinput39);
  xor keyNTinGate_1_7(KeyNOTWire_1[6], keyinput121, keyNTin_Wire_1[7]);
  not KeyNOTGate_1_6(newWire_7, KeyNOTWire_1[6]);
  xnor KeyGate8 (newWire_8, N65, keyinput40);
  xnor KeyGate9 (newWire_9, N89, keyinput41);
  xnor KeyGate10 (newWire_10, N132, keyinput42);
  xor  KeyGate11 (keyNTin_Wire_1[8], N137, keyinput43);
  xor keyNTinGate_1_8(newWire_11, keyinput122, keyNTin_Wire_1[8]);
  xor  KeyGate12 (keyNTin_Wire_1[9], N136, keyinput44);
  xnor keyNTinGate_1_9(newWire_12, keyinput123, keyNTin_Wire_1[9]);
  xnor KeyGate13 (newWire_13, N105, keyinput45);
  xor  KeyGate14 (newWire_14, N97, keyinput46);
  xnor KeyGate15 (newWire_15, N81, keyinput47);
  xnor KeyGate16 (newWire_16, N101, keyinput48);
  xnor KeyGate17 (newWire_17, N5, keyinput49);
  xor  KeyGate18 (keyNTin_Wire_1[10], N37, keyinput50);
  xor keyNTinGate_1_10(newWire_18, keyinput124, keyNTin_Wire_1[10]);
  xor  KeyGate19 (keyNTin_Wire_1[11], N73, keyinput51);
  xnor keyNTinGate_1_11(newWire_19, keyinput125, keyNTin_Wire_1[11]);
  xor  KeyGate20 (keyNTin_Wire_1[12], N1, keyinput52);
  xor keyNTinGate_1_12(KeyNOTWire_1[7], keyinput126, keyNTin_Wire_1[12]);
  not KeyNOTGate_1_7(newWire_20, KeyNOTWire_1[7]);
  xor  KeyGate21 (newWire_21, N13, keyinput53);
  xnor KeyGate22 (newWire_22, N121, keyinput54);
  xor  KeyGate23 (newWire_23, N53, keyinput55);
  xor  KeyGate24 (keyNTin_Wire_1[13], N69, keyinput56);
  xor keyNTinGate_1_13(newWire_24, keyinput127, keyNTin_Wire_1[13]);
  xor  KeyGate25 (keyNTin_Wire_1[14], N113, keyinput57);
  xor keyNTinGate_1_14(KeyNOTWire_1[8], keyinput128, keyNTin_Wire_1[14]);
  not KeyNOTGate_1_8(newWire_25, KeyNOTWire_1[8]);
  xor  KeyGate26 (newWire_26, N33, keyinput58);
  xor  KeyGate27 (newWire_27, N61, keyinput59);
  xor  KeyGate28 (newWire_28, N9, keyinput60);
  xor  KeyGate29 (newWire_29, N41, keyinput61);
  xor  KeyGate30 (newWire_30, N25, keyinput62);
  xor  KeyGate31 (keyNTin_Wire_1[15], N125, keyinput63);
  xor keyNTinGate_1_15(newWire_31, keyinput129, keyNTin_Wire_1[15]);
  xnor KeyGate32 (keyNTin_Wire_1[16], N131, keyinput64);
  xnor keyNTinGate_1_16(KeyNOTWire_1[9], keyinput130, keyNTin_Wire_1[16]);
  not KeyNOTGate_1_9(newWire_32, KeyNOTWire_1[9]);
  xnor KeyGate33 (newWire_33, N135, keyinput65);
  xnor KeyGate34 (keyNTin_Wire_1[17], N117, keyinput66);
  xor keyNTinGate_1_17(KeyNOTWire_1[10], keyinput131, keyNTin_Wire_1[17]);
  not KeyNOTGate_1_10(newWire_34, KeyNOTWire_1[10]);
  xor  KeyGate35 (newWire_35, N85, keyinput67);
  xor  KeyGate36 (keyNTin_Wire_1[18], N57, keyinput68);
  xnor keyNTinGate_1_18(newWire_36, keyinput132, keyNTin_Wire_1[18]);
  xor  KeyGate37 (keyNTin_Wire_1[19], N109, keyinput69);
  xnor keyNTinGate_1_19(KeyNOTWire_1[11], keyinput133, keyNTin_Wire_1[19]);
  not KeyNOTGate_1_11(newWire_37, KeyNOTWire_1[11]);
  xnor KeyGate38 (keyNTin_Wire_1[20], N133, keyinput70);
  xor keyNTinGate_1_20(KeyNOTWire_1[12], keyinput134, keyNTin_Wire_1[20]);
  not KeyNOTGate_1_12(newWire_38, KeyNOTWire_1[12]);
  xnor KeyGate39 (keyNTin_Wire_1[21], N21, keyinput71);
  xnor keyNTinGate_1_21(KeyNOTWire_1[13], keyinput135, keyNTin_Wire_1[21]);
  not KeyNOTGate_1_13(newWire_39, KeyNOTWire_1[13]);
  xor  KeyGate40 (keyNTin_Wire_1[22], N45, keyinput72);
  xor keyNTinGate_1_22(KeyNOTWire_1[14], keyinput136, keyNTin_Wire_1[22]);
  not KeyNOTGate_1_14(newWire_40, KeyNOTWire_1[14]);
  xor  KeyGate41 (newWire_41, N49, keyinput73);
  xor  KeyGate42 (newWire_42, N77, keyinput74);
  xor  KeyGate43 (newWire_43, N17, keyinput75);
  xor  KeyGate44 (newWire_44, N134, keyinput76);
  xnor KeyGate45 (newWire_45, N129, keyinput77);
  xnor KeyGate46 (newWire_46, N130, keyinput78);
  xnor KeyGate47 (keyNTin_Wire_1[23], N29, keyinput79);
  xor keyNTinGate_1_23(newWire_47, keyinput137, keyNTin_Wire_1[23]);
  xnor KeyGate48 (newWire_48, N93, keyinput80);
  xor  KeyGate49 (newWire_49, N65, keyinput81);
  xor  KeyGate50 (newWire_50, N89, keyinput82);
  xor  KeyGate51 (newWire_51, N132, keyinput83);
  xor  KeyGate52 (newWire_52, N137, keyinput84);
  xor  KeyGate53 (keyNTin_Wire_1[24], N136, keyinput85);
  xor keyNTinGate_1_24(newWire_53, keyinput138, keyNTin_Wire_1[24]);
  xor  KeyGate54 (keyNTin_Wire_1[25], N105, keyinput86);
  xnor keyNTinGate_1_25(newWire_54, keyinput139, keyNTin_Wire_1[25]);
  xnor KeyGate55 (newWire_55, N97, keyinput87);
  xnor KeyGate56 (newWire_56, N81, keyinput88);
  xnor KeyGate57 (keyNTin_Wire_1[26], N101, keyinput89);
  xor keyNTinGate_1_26(newWire_57, keyinput140, keyNTin_Wire_1[26]);
  xor  KeyGate58 (keyNTin_Wire_1[27], N5, keyinput90);
  xnor keyNTinGate_1_27(newWire_58, keyinput141, keyNTin_Wire_1[27]);
  xor  KeyGate59 (newWire_59, N37, keyinput91);
  xor  KeyGate60 (newWire_60, N73, keyinput92);
  xor  KeyGate61 (keyNTin_Wire_1[28], N1, keyinput93);
  xnor keyNTinGate_1_28(newWire_61, keyinput142, keyNTin_Wire_1[28]);
  xnor KeyGate62 (keyNTin_Wire_1[29], N13, keyinput94);
  xor keyNTinGate_1_29(KeyNOTWire_1[15], keyinput143, keyNTin_Wire_1[29]);
  not KeyNOTGate_1_15(newWire_62, KeyNOTWire_1[15]);
  xor  KeyGate63 (newWire_63, N121, keyinput95);
  xnor KeyGate64 (newWire_64, N53, keyinput96);
  xor  KeyGate65 (keyNTin_Wire_1[30], N69, keyinput97);
  xor keyNTinGate_1_30(newWire_65, keyinput144, keyNTin_Wire_1[30]);
  xor  KeyGate66 (keyNTin_Wire_1[31], N113, keyinput98);
  xnor keyNTinGate_1_31(KeyNOTWire_1[16], keyinput145, keyNTin_Wire_1[31]);
  not KeyNOTGate_1_16(newWire_66, KeyNOTWire_1[16]);
  xnor KeyGate67 (keyNTin_Wire_1[32], N33, keyinput99);
  xnor keyNTinGate_1_32(KeyNOTWire_1[17], keyinput146, keyNTin_Wire_1[32]);
  not KeyNOTGate_1_17(newWire_67, KeyNOTWire_1[17]);
  xnor KeyGate68 (newWire_68, N61, keyinput100);
  xnor KeyGate69 (keyNTin_Wire_1[33], N9, keyinput101);
  xor keyNTinGate_1_33(KeyNOTWire_1[18], keyinput147, keyNTin_Wire_1[33]);
  not KeyNOTGate_1_18(newWire_69, KeyNOTWire_1[18]);
  xor  KeyGate70 (newWire_70, N41, keyinput102);
  xnor KeyGate71 (newWire_71, N25, keyinput103);
  xor  KeyGate72 (keyNTin_Wire_1[34], N125, keyinput104);
  xor keyNTinGate_1_34(KeyNOTWire_1[19], keyinput148, keyNTin_Wire_1[34]);
  not KeyNOTGate_1_19(newWire_72, KeyNOTWire_1[19]);
  xor  KeyGate73 (newWire_73, N131, keyinput105);
  xnor KeyGate74 (newWire_74, N135, keyinput106);
  xor  KeyGate75 (keyNTin_Wire_1[35], N117, keyinput107);
  xnor keyNTinGate_1_35(newWire_75, keyinput149, keyNTin_Wire_1[35]);
  xnor KeyGate76 (newWire_76, N85, keyinput108);
  xor  KeyGate77 (keyNTin_Wire_1[36], N57, keyinput109);
  xor keyNTinGate_1_36(newWire_77, keyinput150, keyNTin_Wire_1[36]);
  xor  KeyGate78 (newWire_78, N109, keyinput110);
  xnor KeyGate79 (keyNTin_Wire_1[37], N133, keyinput111);
  xnor keyNTinGate_1_37(KeyNOTWire_1[20], keyinput151, keyNTin_Wire_1[37]);
  not KeyNOTGate_1_20(newWire_79, KeyNOTWire_1[20]);
  xor  KeyGate80 (newWire_80, N21, keyinput112);
  xnor KeyGate81 (keyNTin_Wire_1[38], N45, keyinput113);
  xnor keyNTinGate_1_38(newWire_81, keyinput152, keyNTin_Wire_1[38]);
  and some_function (keyNTin_Wire_1[39], newWire_0, newWire_1, newWire_2, newWire_3, newWire_4, newWire_5, newWire_6, newWire_7, newWire_8, newWire_9, newWire_10, newWire_11, newWire_12, newWire_13, newWire_14, newWire_15, newWire_16, newWire_17, newWire_18, newWire_19, newWire_20, newWire_21, newWire_22, newWire_23, newWire_24, newWire_25, newWire_26, newWire_27, newWire_28, newWire_29, newWire_30, newWire_31, newWire_32, newWire_33, newWire_34, newWire_35, newWire_36, newWire_37, newWire_38, newWire_39, newWire_40 );
  xnor keyNTinGate_1_39(KeyNOTWire_1[21], keyinput153, keyNTin_Wire_1[39]);
  not KeyNOTGate_1_21(newWire_82, KeyNOTWire_1[21]);
  nand compl_function (newWire_83, newWire_41, newWire_42, newWire_43, newWire_44, newWire_45, newWire_46, newWire_47, newWire_48, newWire_49, newWire_50, newWire_51, newWire_52, newWire_53, newWire_54, newWire_55, newWire_56, newWire_57, newWire_58, newWire_59, newWire_60, newWire_61, newWire_62, newWire_63, newWire_64, newWire_65, newWire_66, newWire_67, newWire_68, newWire_69, newWire_70, newWire_71, newWire_72, newWire_73, newWire_74, newWire_75, newWire_76, newWire_77, newWire_78, newWire_79, newWire_80, newWire_81);
  and finalAND (keyNTin_Wire_1[40], newWire_82, newWire_83);
  xnor keyNTinGate_1_40(KeyWire_0_2, keyinput154, keyNTin_Wire_1[40]);

endmodule /* AntiSAT */
