`timescale 1ns / 1ps
// Verilog
// c880
// Ninputs 60
// Noutputs 26
// NtotalGates 383
// NAND4 13
// AND3 12
// NAND2 60
// NAND3 14
// AND2 105
// OR2 29
// NOT1 63
// NOR2 61
// BUFF1 26

module top (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
                  N865,N866,N874,N878,N879,N880,
        keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4,
        keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9,
        keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14,
        keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19,
        keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24,
        keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29,
        keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34,
        keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39,
        keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44,
        keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49,
        keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54,
        keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59,
        keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64,
        keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69,
        keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74,
        keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79,
        keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84,
        keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89,
        keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94,
        keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99,
        keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104,
        keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109,
        keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114,
        keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119,
        keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124,
        keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129,
        keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134,
        keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139,
        keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144,
        keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149,
        keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154,
        keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159,
        keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164,
        keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169,
        keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174,
        keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179,
        keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184,
        keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189,
        keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194,
        keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199,
        keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204,
        keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209,
        keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214,
        keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219,
        keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224,
        keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229,
        keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234,
        keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239,
        keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244,
        keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249,
        keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254,
        keyIn_0_255);

  input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4;
  input keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9;
  input keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14;
  input keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19;
  input keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24;
  input keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29;
  input keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34;
  input keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39;
  input keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44;
  input keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49;
  input keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54;
  input keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59;
  input keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64;
  input keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69;
  input keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74;
  input keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79;
  input keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84;
  input keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89;
  input keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94;
  input keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99;
  input keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104;
  input keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109;
  input keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114;
  input keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119;
  input keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124;
  input keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129;
  input keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134;
  input keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139;
  input keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144;
  input keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149;
  input keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154;
  input keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159;
  input keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164;
  input keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169;
  input keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174;
  input keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179;
  input keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184;
  input keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189;
  input keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194;
  input keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199;
  input keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204;
  input keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209;
  input keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214;
  input keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219;
  input keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224;
  input keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229;
  input keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234;
  input keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239;
  input keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244;
  input keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249;
  input keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254;
  input keyIn_0_255;

  wire [0:255] KeyWire_0;
  wire [0:125] KeyNOTWire_0;

input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;

output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;

wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877;

nand NAND4_1 (N269, N1, N8, N13, N17);
nand NAND4_2 (N270, N1, N26, N13, N17);
and AND3_3 (N273, N29, N36, N42);
  and AND3_4 (KeyWire_0[0], N1, N26, N51);
  xnor KeyGate_0_0(KeyNOTWire_0[0], keyIn_0_0, KeyWire_0[0]);
  not KeyNOTGate_0_0(N276, KeyNOTWire_0[0]);
  nand NAND4_5 (KeyWire_0[1], N1, N8, N51, N17);
  xnor KeyGate_0_1(N279, keyIn_0_1, KeyWire_0[1]);
  nand NAND4_6 (KeyWire_0[2], N1, N8, N13, N55);
  xor KeyGate_0_2(N280, keyIn_0_2, KeyWire_0[2]);
  nand NAND4_7 (KeyWire_0[3], N59, N42, N68, N72);
  xor KeyGate_0_3(N284, keyIn_0_3, KeyWire_0[3]);
nand NAND2_8 (N285, N29, N68);
nand NAND3_9 (N286, N59, N68, N74);
  and AND3_10 (KeyWire_0[4], N29, N75, N80);
  xnor KeyGate_0_4(N287, keyIn_0_4, KeyWire_0[4]);
and AND3_11 (N290, N29, N75, N42);
and AND3_12 (N291, N29, N36, N80);
and AND3_13 (N292, N29, N36, N42);
and AND3_14 (N293, N59, N75, N80);
  and AND3_15 (KeyWire_0[5], N59, N75, N42);
  xnor KeyGate_0_5(N294, keyIn_0_5, KeyWire_0[5]);
and AND3_16 (N295, N59, N36, N80);
and AND3_17 (N296, N59, N36, N42);
and AND2_18 (N297, N85, N86);
or OR2_19 (N298, N87, N88);
nand NAND2_20 (N301, N91, N96);
or OR2_21 (N302, N91, N96);
nand NAND2_22 (N303, N101, N106);
or OR2_23 (N304, N101, N106);
  nand NAND2_24 (KeyWire_0[6], N111, N116);
  xnor KeyGate_0_6(KeyNOTWire_0[1], keyIn_0_6, KeyWire_0[6]);
  not KeyNOTGate_0_1(N305, KeyNOTWire_0[1]);
or OR2_25 (N306, N111, N116);
nand NAND2_26 (N307, N121, N126);
or OR2_27 (N308, N121, N126);
  and AND2_28 (KeyWire_0[7], N8, N138);
  xor KeyGate_0_7(KeyNOTWire_0[2], keyIn_0_7, KeyWire_0[7]);
  not KeyNOTGate_0_2(N309, KeyNOTWire_0[2]);
  not NOT1_29 (KeyWire_0[8], N268);
  xnor KeyGate_0_8(KeyNOTWire_0[3], keyIn_0_8, KeyWire_0[8]);
  not KeyNOTGate_0_3(N310, KeyNOTWire_0[3]);
  and AND2_30 (KeyWire_0[9], N51, N138);
  xnor KeyGate_0_9(KeyNOTWire_0[4], keyIn_0_9, KeyWire_0[9]);
  not KeyNOTGate_0_4(N316, KeyNOTWire_0[4]);
  and AND2_31 (KeyWire_0[10], N17, N138);
  xor KeyGate_0_10(KeyNOTWire_0[5], keyIn_0_10, KeyWire_0[10]);
  not KeyNOTGate_0_5(N317, KeyNOTWire_0[5]);
  and AND2_32 (KeyWire_0[11], N152, N138);
  xnor KeyGate_0_11(N318, keyIn_0_11, KeyWire_0[11]);
  nand NAND2_33 (KeyWire_0[12], N59, N156);
  xnor KeyGate_0_12(KeyNOTWire_0[6], keyIn_0_12, KeyWire_0[12]);
  not KeyNOTGate_0_6(N319, KeyNOTWire_0[6]);
  nor NOR2_34 (KeyWire_0[13], N17, N42);
  xor KeyGate_0_13(N322, keyIn_0_13, KeyWire_0[13]);
  and AND2_35 (KeyWire_0[14], N17, N42);
  xor KeyGate_0_14(N323, keyIn_0_14, KeyWire_0[14]);
nand NAND2_36 (N324, N159, N165);
or OR2_37 (N325, N159, N165);
nand NAND2_38 (N326, N171, N177);
or OR2_39 (N327, N171, N177);
nand NAND2_40 (N328, N183, N189);
or OR2_41 (N329, N183, N189);
nand NAND2_42 (N330, N195, N201);
or OR2_43 (N331, N195, N201);
  and AND2_44 (KeyWire_0[15], N210, N91);
  xnor KeyGate_0_15(KeyNOTWire_0[7], keyIn_0_15, KeyWire_0[15]);
  not KeyNOTGate_0_7(N332, KeyNOTWire_0[7]);
and AND2_45 (N333, N210, N96);
and AND2_46 (N334, N210, N101);
and AND2_47 (N335, N210, N106);
  and AND2_48 (KeyWire_0[16], N210, N111);
  xnor KeyGate_0_16(N336, keyIn_0_16, KeyWire_0[16]);
and AND2_49 (N337, N255, N259);
and AND2_50 (N338, N210, N116);
and AND2_51 (N339, N255, N260);
  and AND2_52 (KeyWire_0[17], N210, N121);
  xor KeyGate_0_17(N340, keyIn_0_17, KeyWire_0[17]);
and AND2_53 (N341, N255, N267);
not NOT1_54 (N342, N269);
not NOT1_55 (N343, N273);
or OR2_56 (N344, N270, N273);
  not NOT1_57 (KeyWire_0[18], N276);
  xnor KeyGate_0_18(KeyNOTWire_0[8], keyIn_0_18, KeyWire_0[18]);
  not KeyNOTGate_0_8(N345, KeyNOTWire_0[8]);
not NOT1_58 (N346, N276);
  not NOT1_59 (KeyWire_0[19], N279);
  xor KeyGate_0_19(KeyNOTWire_0[9], keyIn_0_19, KeyWire_0[19]);
  not KeyNOTGate_0_9(N347, KeyNOTWire_0[9]);
  nor NOR2_60 (KeyWire_0[20], N280, N284);
  xor KeyGate_0_20(N348, keyIn_0_20, KeyWire_0[20]);
or OR2_61 (N349, N280, N285);
or OR2_62 (N350, N280, N286);
not NOT1_63 (N351, N293);
  not NOT1_64 (KeyWire_0[21], N294);
  xor KeyGate_0_21(KeyNOTWire_0[10], keyIn_0_21, KeyWire_0[21]);
  not KeyNOTGate_0_10(N352, KeyNOTWire_0[10]);
not NOT1_65 (N353, N295);
not NOT1_66 (N354, N296);
nand NAND2_67 (N355, N89, N298);
  and AND2_68 (KeyWire_0[22], N90, N298);
  xnor KeyGate_0_22(N356, keyIn_0_22, KeyWire_0[22]);
nand NAND2_69 (N357, N301, N302);
nand NAND2_70 (N360, N303, N304);
nand NAND2_71 (N363, N305, N306);
nand NAND2_72 (N366, N307, N308);
  not NOT1_73 (KeyWire_0[23], N310);
  xor KeyGate_0_23(N369, keyIn_0_23, KeyWire_0[23]);
  nor NOR2_74 (KeyWire_0[24], N322, N323);
  xor KeyGate_0_24(N375, keyIn_0_24, KeyWire_0[24]);
nand NAND2_75 (N376, N324, N325);
nand NAND2_76 (N379, N326, N327);
nand NAND2_77 (N382, N328, N329);
nand NAND2_78 (N385, N330, N331);
buf BUFF1_79 (N388, N290);
buf BUFF1_80 (N389, N291);
buf BUFF1_81 (N390, N292);
buf BUFF1_82 (N391, N297);
or OR2_83 (N392, N270, N343);
  not NOT1_84 (KeyWire_0[25], N345);
  xor KeyGate_0_25(KeyNOTWire_0[11], keyIn_0_25, KeyWire_0[25]);
  not KeyNOTGate_0_11(N393, KeyNOTWire_0[11]);
  not NOT1_85 (KeyWire_0[26], N346);
  xor KeyGate_0_26(KeyNOTWire_0[12], keyIn_0_26, KeyWire_0[26]);
  not KeyNOTGate_0_12(N399, KeyNOTWire_0[12]);
  and AND2_86 (KeyWire_0[27], N348, N73);
  xnor KeyGate_0_27(KeyNOTWire_0[13], keyIn_0_27, KeyWire_0[27]);
  not KeyNOTGate_0_13(N400, KeyNOTWire_0[13]);
not NOT1_87 (N401, N349);
not NOT1_88 (N402, N350);
not NOT1_89 (N403, N355);
not NOT1_90 (N404, N357);
not NOT1_91 (N405, N360);
and AND2_92 (N406, N357, N360);
not NOT1_93 (N407, N363);
not NOT1_94 (N408, N366);
and AND2_95 (N409, N363, N366);
  nand NAND2_96 (KeyWire_0[28], N347, N352);
  xor KeyGate_0_28(KeyNOTWire_0[14], keyIn_0_28, KeyWire_0[28]);
  not KeyNOTGate_0_14(N410, KeyNOTWire_0[14]);
not NOT1_97 (N411, N376);
not NOT1_98 (N412, N379);
and AND2_99 (N413, N376, N379);
not NOT1_100 (N414, N382);
not NOT1_101 (N415, N385);
and AND2_102 (N416, N382, N385);
  and AND2_103 (KeyWire_0[29], N210, N369);
  xor KeyGate_0_29(N417, keyIn_0_29, KeyWire_0[29]);
buf BUFF1_104 (N418, N342);
buf BUFF1_105 (N419, N344);
buf BUFF1_106 (N420, N351);
buf BUFF1_107 (N421, N353);
buf BUFF1_108 (N422, N354);
buf BUFF1_109 (N423, N356);
  not NOT1_110 (KeyWire_0[30], N400);
  xor KeyGate_0_30(N424, keyIn_0_30, KeyWire_0[30]);
and AND2_111 (N425, N404, N405);
and AND2_112 (N426, N407, N408);
  and AND3_113 (KeyWire_0[31], N319, N393, N55);
  xor KeyGate_0_31(KeyNOTWire_0[15], keyIn_0_31, KeyWire_0[31]);
  not KeyNOTGate_0_15(N427, KeyNOTWire_0[15]);
  and AND3_114 (KeyWire_0[32], N393, N17, N287);
  xnor KeyGate_0_32(N432, keyIn_0_32, KeyWire_0[32]);
  nand NAND3_115 (KeyWire_0[33], N393, N287, N55);
  xnor KeyGate_0_33(N437, keyIn_0_33, KeyWire_0[33]);
  nand NAND4_116 (KeyWire_0[34], N375, N59, N156, N393);
  xor KeyGate_0_34(KeyNOTWire_0[16], keyIn_0_34, KeyWire_0[34]);
  not KeyNOTGate_0_16(N442, KeyNOTWire_0[16]);
  nand NAND3_117 (KeyWire_0[35], N393, N319, N17);
  xor KeyGate_0_35(KeyNOTWire_0[17], keyIn_0_35, KeyWire_0[35]);
  not KeyNOTGate_0_17(N443, KeyNOTWire_0[17]);
and AND2_118 (N444, N411, N412);
and AND2_119 (N445, N414, N415);
buf BUFF1_120 (N446, N392);
buf BUFF1_121 (N447, N399);
buf BUFF1_122 (N448, N401);
buf BUFF1_123 (N449, N402);
buf BUFF1_124 (N450, N403);
  not NOT1_125 (KeyWire_0[36], N424);
  xnor KeyGate_0_36(N451, keyIn_0_36, KeyWire_0[36]);
nor NOR2_126 (N460, N406, N425);
nor NOR2_127 (N463, N409, N426);
  nand NAND2_128 (KeyWire_0[37], N442, N410);
  xnor KeyGate_0_37(N466, keyIn_0_37, KeyWire_0[37]);
  and AND2_129 (KeyWire_0[38], N143, N427);
  xnor KeyGate_0_38(N475, keyIn_0_38, KeyWire_0[38]);
  and AND2_130 (KeyWire_0[39], N310, N432);
  xor KeyGate_0_39(N476, keyIn_0_39, KeyWire_0[39]);
  and AND2_131 (KeyWire_0[40], N146, N427);
  xor KeyGate_0_40(N477, keyIn_0_40, KeyWire_0[40]);
  and AND2_132 (KeyWire_0[41], N310, N432);
  xor KeyGate_0_41(KeyNOTWire_0[18], keyIn_0_41, KeyWire_0[41]);
  not KeyNOTGate_0_18(N478, KeyNOTWire_0[18]);
  and AND2_133 (KeyWire_0[42], N149, N427);
  xor KeyGate_0_42(N479, keyIn_0_42, KeyWire_0[42]);
  and AND2_134 (KeyWire_0[43], N310, N432);
  xor KeyGate_0_43(KeyNOTWire_0[19], keyIn_0_43, KeyWire_0[43]);
  not KeyNOTGate_0_19(N480, KeyNOTWire_0[19]);
  and AND2_135 (KeyWire_0[44], N153, N427);
  xnor KeyGate_0_44(N481, keyIn_0_44, KeyWire_0[44]);
  and AND2_136 (KeyWire_0[45], N310, N432);
  xnor KeyGate_0_45(KeyNOTWire_0[20], keyIn_0_45, KeyWire_0[45]);
  not KeyNOTGate_0_20(N482, KeyNOTWire_0[20]);
  nand NAND2_137 (KeyWire_0[46], N443, N1);
  xnor KeyGate_0_46(N483, keyIn_0_46, KeyWire_0[46]);
  or OR2_138 (KeyWire_0[47], N369, N437);
  xnor KeyGate_0_47(N488, keyIn_0_47, KeyWire_0[47]);
  or OR2_139 (KeyWire_0[48], N369, N437);
  xnor KeyGate_0_48(KeyNOTWire_0[21], keyIn_0_48, KeyWire_0[48]);
  not KeyNOTGate_0_21(N489, KeyNOTWire_0[21]);
  or OR2_140 (KeyWire_0[49], N369, N437);
  xor KeyGate_0_49(KeyNOTWire_0[22], keyIn_0_49, KeyWire_0[49]);
  not KeyNOTGate_0_22(N490, KeyNOTWire_0[22]);
  or OR2_141 (KeyWire_0[50], N369, N437);
  xnor KeyGate_0_50(KeyNOTWire_0[23], keyIn_0_50, KeyWire_0[50]);
  not KeyNOTGate_0_23(N491, KeyNOTWire_0[23]);
nor NOR2_142 (N492, N413, N444);
nor NOR2_143 (N495, N416, N445);
nand NAND2_144 (N498, N130, N460);
or OR2_145 (N499, N130, N460);
nand NAND2_146 (N500, N463, N135);
or OR2_147 (N501, N463, N135);
  and AND2_148 (KeyWire_0[51], N91, N466);
  xnor KeyGate_0_51(KeyNOTWire_0[24], keyIn_0_51, KeyWire_0[51]);
  not KeyNOTGate_0_24(N502, KeyNOTWire_0[24]);
  nor NOR2_149 (KeyWire_0[52], N475, N476);
  xor KeyGate_0_52(N503, keyIn_0_52, KeyWire_0[52]);
  and AND2_150 (KeyWire_0[53], N96, N466);
  xnor KeyGate_0_53(N504, keyIn_0_53, KeyWire_0[53]);
  nor NOR2_151 (KeyWire_0[54], N477, N478);
  xor KeyGate_0_54(KeyNOTWire_0[25], keyIn_0_54, KeyWire_0[54]);
  not KeyNOTGate_0_25(N505, KeyNOTWire_0[25]);
  and AND2_152 (KeyWire_0[55], N101, N466);
  xnor KeyGate_0_55(N506, keyIn_0_55, KeyWire_0[55]);
  nor NOR2_153 (KeyWire_0[56], N479, N480);
  xor KeyGate_0_56(N507, keyIn_0_56, KeyWire_0[56]);
  and AND2_154 (KeyWire_0[57], N106, N466);
  xnor KeyGate_0_57(KeyNOTWire_0[26], keyIn_0_57, KeyWire_0[57]);
  not KeyNOTGate_0_26(N508, KeyNOTWire_0[26]);
  nor NOR2_155 (KeyWire_0[58], N481, N482);
  xnor KeyGate_0_58(KeyNOTWire_0[27], keyIn_0_58, KeyWire_0[58]);
  not KeyNOTGate_0_27(N509, KeyNOTWire_0[27]);
  and AND2_156 (KeyWire_0[59], N143, N483);
  xor KeyGate_0_59(N510, keyIn_0_59, KeyWire_0[59]);
  and AND2_157 (KeyWire_0[60], N111, N466);
  xnor KeyGate_0_60(N511, keyIn_0_60, KeyWire_0[60]);
  and AND2_158 (KeyWire_0[61], N146, N483);
  xor KeyGate_0_61(N512, keyIn_0_61, KeyWire_0[61]);
  and AND2_159 (KeyWire_0[62], N116, N466);
  xor KeyGate_0_62(KeyNOTWire_0[28], keyIn_0_62, KeyWire_0[62]);
  not KeyNOTGate_0_28(N513, KeyNOTWire_0[28]);
  and AND2_160 (KeyWire_0[63], N149, N483);
  xnor KeyGate_0_63(N514, keyIn_0_63, KeyWire_0[63]);
  and AND2_161 (KeyWire_0[64], N121, N466);
  xnor KeyGate_0_64(N515, keyIn_0_64, KeyWire_0[64]);
  and AND2_162 (KeyWire_0[65], N153, N483);
  xnor KeyGate_0_65(KeyNOTWire_0[29], keyIn_0_65, KeyWire_0[65]);
  not KeyNOTGate_0_29(N516, KeyNOTWire_0[29]);
  and AND2_163 (KeyWire_0[66], N126, N466);
  xor KeyGate_0_66(N517, keyIn_0_66, KeyWire_0[66]);
nand NAND2_164 (N518, N130, N492);
or OR2_165 (N519, N130, N492);
nand NAND2_166 (N520, N495, N207);
or OR2_167 (N521, N495, N207);
  and AND2_168 (KeyWire_0[67], N451, N159);
  xor KeyGate_0_67(KeyNOTWire_0[30], keyIn_0_67, KeyWire_0[67]);
  not KeyNOTGate_0_30(N522, KeyNOTWire_0[30]);
  and AND2_169 (KeyWire_0[68], N451, N165);
  xor KeyGate_0_68(KeyNOTWire_0[31], keyIn_0_68, KeyWire_0[68]);
  not KeyNOTGate_0_31(N523, KeyNOTWire_0[31]);
  and AND2_170 (KeyWire_0[69], N451, N171);
  xor KeyGate_0_69(KeyNOTWire_0[32], keyIn_0_69, KeyWire_0[69]);
  not KeyNOTGate_0_32(N524, KeyNOTWire_0[32]);
  and AND2_171 (KeyWire_0[70], N451, N177);
  xor KeyGate_0_70(N525, keyIn_0_70, KeyWire_0[70]);
  and AND2_172 (KeyWire_0[71], N451, N183);
  xor KeyGate_0_71(N526, keyIn_0_71, KeyWire_0[71]);
  nand NAND2_173 (KeyWire_0[72], N451, N189);
  xor KeyGate_0_72(N527, keyIn_0_72, KeyWire_0[72]);
nand NAND2_174 (N528, N451, N195);
nand NAND2_175 (N529, N451, N201);
nand NAND2_176 (N530, N498, N499);
nand NAND2_177 (N533, N500, N501);
  nor NOR2_178 (KeyWire_0[73], N309, N502);
  xor KeyGate_0_73(KeyNOTWire_0[33], keyIn_0_73, KeyWire_0[73]);
  not KeyNOTGate_0_33(N536, KeyNOTWire_0[33]);
  nor NOR2_179 (KeyWire_0[74], N316, N504);
  xor KeyGate_0_74(KeyNOTWire_0[34], keyIn_0_74, KeyWire_0[74]);
  not KeyNOTGate_0_34(N537, KeyNOTWire_0[34]);
  nor NOR2_180 (KeyWire_0[75], N317, N506);
  xnor KeyGate_0_75(N538, keyIn_0_75, KeyWire_0[75]);
  nor NOR2_181 (KeyWire_0[76], N318, N508);
  xnor KeyGate_0_76(N539, keyIn_0_76, KeyWire_0[76]);
  nor NOR2_182 (KeyWire_0[77], N510, N511);
  xor KeyGate_0_77(KeyNOTWire_0[35], keyIn_0_77, KeyWire_0[77]);
  not KeyNOTGate_0_35(N540, KeyNOTWire_0[35]);
  nor NOR2_183 (KeyWire_0[78], N512, N513);
  xnor KeyGate_0_78(KeyNOTWire_0[36], keyIn_0_78, KeyWire_0[78]);
  not KeyNOTGate_0_36(N541, KeyNOTWire_0[36]);
  nor NOR2_184 (KeyWire_0[79], N514, N515);
  xor KeyGate_0_79(KeyNOTWire_0[37], keyIn_0_79, KeyWire_0[79]);
  not KeyNOTGate_0_37(N542, KeyNOTWire_0[37]);
  nor NOR2_185 (KeyWire_0[80], N516, N517);
  xor KeyGate_0_80(KeyNOTWire_0[38], keyIn_0_80, KeyWire_0[80]);
  not KeyNOTGate_0_38(N543, KeyNOTWire_0[38]);
nand NAND2_186 (N544, N518, N519);
nand NAND2_187 (N547, N520, N521);
not NOT1_188 (N550, N530);
not NOT1_189 (N551, N533);
and AND2_190 (N552, N530, N533);
  nand NAND2_191 (KeyWire_0[81], N536, N503);
  xnor KeyGate_0_81(KeyNOTWire_0[39], keyIn_0_81, KeyWire_0[81]);
  not KeyNOTGate_0_39(N553, KeyNOTWire_0[39]);
  nand NAND2_192 (KeyWire_0[82], N537, N505);
  xnor KeyGate_0_82(N557, keyIn_0_82, KeyWire_0[82]);
  nand NAND2_193 (KeyWire_0[83], N538, N507);
  xor KeyGate_0_83(KeyNOTWire_0[40], keyIn_0_83, KeyWire_0[83]);
  not KeyNOTGate_0_40(N561, KeyNOTWire_0[40]);
  nand NAND2_194 (KeyWire_0[84], N539, N509);
  xnor KeyGate_0_84(N565, keyIn_0_84, KeyWire_0[84]);
  nand NAND2_195 (KeyWire_0[85], N488, N540);
  xor KeyGate_0_85(KeyNOTWire_0[41], keyIn_0_85, KeyWire_0[85]);
  not KeyNOTGate_0_41(N569, KeyNOTWire_0[41]);
  nand NAND2_196 (KeyWire_0[86], N489, N541);
  xnor KeyGate_0_86(KeyNOTWire_0[42], keyIn_0_86, KeyWire_0[86]);
  not KeyNOTGate_0_42(N573, KeyNOTWire_0[42]);
  nand NAND2_197 (KeyWire_0[87], N490, N542);
  xor KeyGate_0_87(KeyNOTWire_0[43], keyIn_0_87, KeyWire_0[87]);
  not KeyNOTGate_0_43(N577, KeyNOTWire_0[43]);
  nand NAND2_198 (KeyWire_0[88], N491, N543);
  xnor KeyGate_0_88(N581, keyIn_0_88, KeyWire_0[88]);
not NOT1_199 (N585, N544);
not NOT1_200 (N586, N547);
and AND2_201 (N587, N544, N547);
and AND2_202 (N588, N550, N551);
and AND2_203 (N589, N585, N586);
  nand NAND2_204 (KeyWire_0[89], N553, N159);
  xnor KeyGate_0_89(KeyNOTWire_0[44], keyIn_0_89, KeyWire_0[89]);
  not KeyNOTGate_0_44(N590, KeyNOTWire_0[44]);
  or OR2_205 (KeyWire_0[90], N553, N159);
  xor KeyGate_0_90(N593, keyIn_0_90, KeyWire_0[90]);
  and AND2_206 (KeyWire_0[91], N246, N553);
  xor KeyGate_0_91(N596, keyIn_0_91, KeyWire_0[91]);
  nand NAND2_207 (KeyWire_0[92], N557, N165);
  xor KeyGate_0_92(N597, keyIn_0_92, KeyWire_0[92]);
  or OR2_208 (KeyWire_0[93], N557, N165);
  xor KeyGate_0_93(N600, keyIn_0_93, KeyWire_0[93]);
  and AND2_209 (KeyWire_0[94], N246, N557);
  xor KeyGate_0_94(KeyNOTWire_0[45], keyIn_0_94, KeyWire_0[94]);
  not KeyNOTGate_0_45(N605, KeyNOTWire_0[45]);
  nand NAND2_210 (KeyWire_0[95], N561, N171);
  xor KeyGate_0_95(N606, keyIn_0_95, KeyWire_0[95]);
  or OR2_211 (KeyWire_0[96], N561, N171);
  xnor KeyGate_0_96(N609, keyIn_0_96, KeyWire_0[96]);
  and AND2_212 (KeyWire_0[97], N246, N561);
  xor KeyGate_0_97(N615, keyIn_0_97, KeyWire_0[97]);
  nand NAND2_213 (KeyWire_0[98], N565, N177);
  xor KeyGate_0_98(KeyNOTWire_0[46], keyIn_0_98, KeyWire_0[98]);
  not KeyNOTGate_0_46(N616, KeyNOTWire_0[46]);
  or OR2_214 (KeyWire_0[99], N565, N177);
  xnor KeyGate_0_99(KeyNOTWire_0[47], keyIn_0_99, KeyWire_0[99]);
  not KeyNOTGate_0_47(N619, KeyNOTWire_0[47]);
  and AND2_215 (KeyWire_0[100], N246, N565);
  xor KeyGate_0_100(N624, keyIn_0_100, KeyWire_0[100]);
  nand NAND2_216 (KeyWire_0[101], N569, N183);
  xor KeyGate_0_101(KeyNOTWire_0[48], keyIn_0_101, KeyWire_0[101]);
  not KeyNOTGate_0_48(N625, KeyNOTWire_0[48]);
  or OR2_217 (KeyWire_0[102], N569, N183);
  xor KeyGate_0_102(N628, keyIn_0_102, KeyWire_0[102]);
  and AND2_218 (KeyWire_0[103], N246, N569);
  xor KeyGate_0_103(N631, keyIn_0_103, KeyWire_0[103]);
  nand NAND2_219 (KeyWire_0[104], N573, N189);
  xnor KeyGate_0_104(N632, keyIn_0_104, KeyWire_0[104]);
  or OR2_220 (KeyWire_0[105], N573, N189);
  xnor KeyGate_0_105(N635, keyIn_0_105, KeyWire_0[105]);
  and AND2_221 (KeyWire_0[106], N246, N573);
  xnor KeyGate_0_106(N640, keyIn_0_106, KeyWire_0[106]);
  nand NAND2_222 (KeyWire_0[107], N577, N195);
  xor KeyGate_0_107(KeyNOTWire_0[49], keyIn_0_107, KeyWire_0[107]);
  not KeyNOTGate_0_49(N641, KeyNOTWire_0[49]);
  or OR2_223 (KeyWire_0[108], N577, N195);
  xor KeyGate_0_108(KeyNOTWire_0[50], keyIn_0_108, KeyWire_0[108]);
  not KeyNOTGate_0_50(N644, KeyNOTWire_0[50]);
  and AND2_224 (KeyWire_0[109], N246, N577);
  xnor KeyGate_0_109(KeyNOTWire_0[51], keyIn_0_109, KeyWire_0[109]);
  not KeyNOTGate_0_51(N650, KeyNOTWire_0[51]);
  nand NAND2_225 (KeyWire_0[110], N581, N201);
  xnor KeyGate_0_110(N651, keyIn_0_110, KeyWire_0[110]);
  or OR2_226 (KeyWire_0[111], N581, N201);
  xor KeyGate_0_111(KeyNOTWire_0[52], keyIn_0_111, KeyWire_0[111]);
  not KeyNOTGate_0_52(N654, KeyNOTWire_0[52]);
  and AND2_227 (KeyWire_0[112], N246, N581);
  xor KeyGate_0_112(KeyNOTWire_0[53], keyIn_0_112, KeyWire_0[112]);
  not KeyNOTGate_0_53(N659, KeyNOTWire_0[53]);
nor NOR2_228 (N660, N552, N588);
nor NOR2_229 (N661, N587, N589);
  not NOT1_230 (KeyWire_0[113], N590);
  xor KeyGate_0_113(N662, keyIn_0_113, KeyWire_0[113]);
  and AND2_231 (KeyWire_0[114], N593, N590);
  xnor KeyGate_0_114(N665, keyIn_0_114, KeyWire_0[114]);
  nor NOR2_232 (KeyWire_0[115], N596, N522);
  xor KeyGate_0_115(N669, keyIn_0_115, KeyWire_0[115]);
  not NOT1_233 (KeyWire_0[116], N597);
  xor KeyGate_0_116(N670, keyIn_0_116, KeyWire_0[116]);
  and AND2_234 (KeyWire_0[117], N600, N597);
  xnor KeyGate_0_117(KeyNOTWire_0[54], keyIn_0_117, KeyWire_0[117]);
  not KeyNOTGate_0_54(N673, KeyNOTWire_0[54]);
  nor NOR2_235 (KeyWire_0[118], N605, N523);
  xor KeyGate_0_118(KeyNOTWire_0[55], keyIn_0_118, KeyWire_0[118]);
  not KeyNOTGate_0_55(N677, KeyNOTWire_0[55]);
  not NOT1_236 (KeyWire_0[119], N606);
  xor KeyGate_0_119(KeyNOTWire_0[56], keyIn_0_119, KeyWire_0[119]);
  not KeyNOTGate_0_56(N678, KeyNOTWire_0[56]);
  and AND2_237 (KeyWire_0[120], N609, N606);
  xnor KeyGate_0_120(KeyNOTWire_0[57], keyIn_0_120, KeyWire_0[120]);
  not KeyNOTGate_0_57(N682, KeyNOTWire_0[57]);
  nor NOR2_238 (KeyWire_0[121], N615, N524);
  xnor KeyGate_0_121(KeyNOTWire_0[58], keyIn_0_121, KeyWire_0[121]);
  not KeyNOTGate_0_58(N686, KeyNOTWire_0[58]);
  not NOT1_239 (KeyWire_0[122], N616);
  xor KeyGate_0_122(KeyNOTWire_0[59], keyIn_0_122, KeyWire_0[122]);
  not KeyNOTGate_0_59(N687, KeyNOTWire_0[59]);
  and AND2_240 (KeyWire_0[123], N619, N616);
  xnor KeyGate_0_123(KeyNOTWire_0[60], keyIn_0_123, KeyWire_0[123]);
  not KeyNOTGate_0_60(N692, KeyNOTWire_0[60]);
  nor NOR2_241 (KeyWire_0[124], N624, N525);
  xnor KeyGate_0_124(N696, keyIn_0_124, KeyWire_0[124]);
  not NOT1_242 (KeyWire_0[125], N625);
  xnor KeyGate_0_125(KeyNOTWire_0[61], keyIn_0_125, KeyWire_0[125]);
  not KeyNOTGate_0_61(N697, KeyNOTWire_0[61]);
  and AND2_243 (KeyWire_0[126], N628, N625);
  xor KeyGate_0_126(N700, keyIn_0_126, KeyWire_0[126]);
  nor NOR2_244 (KeyWire_0[127], N631, N526);
  xor KeyGate_0_127(N704, keyIn_0_127, KeyWire_0[127]);
  not NOT1_245 (KeyWire_0[128], N632);
  xor KeyGate_0_128(N705, keyIn_0_128, KeyWire_0[128]);
  and AND2_246 (KeyWire_0[129], N635, N632);
  xnor KeyGate_0_129(KeyNOTWire_0[62], keyIn_0_129, KeyWire_0[129]);
  not KeyNOTGate_0_62(N708, KeyNOTWire_0[62]);
  nor NOR2_247 (KeyWire_0[130], N337, N640);
  xor KeyGate_0_130(KeyNOTWire_0[63], keyIn_0_130, KeyWire_0[130]);
  not KeyNOTGate_0_63(N712, KeyNOTWire_0[63]);
  not NOT1_248 (KeyWire_0[131], N641);
  xnor KeyGate_0_131(KeyNOTWire_0[64], keyIn_0_131, KeyWire_0[131]);
  not KeyNOTGate_0_64(N713, KeyNOTWire_0[64]);
  and AND2_249 (KeyWire_0[132], N644, N641);
  xor KeyGate_0_132(N717, keyIn_0_132, KeyWire_0[132]);
  nor NOR2_250 (KeyWire_0[133], N339, N650);
  xnor KeyGate_0_133(N721, keyIn_0_133, KeyWire_0[133]);
  not NOT1_251 (KeyWire_0[134], N651);
  xnor KeyGate_0_134(N722, keyIn_0_134, KeyWire_0[134]);
  and AND2_252 (KeyWire_0[135], N654, N651);
  xor KeyGate_0_135(KeyNOTWire_0[65], keyIn_0_135, KeyWire_0[135]);
  not KeyNOTGate_0_65(N727, KeyNOTWire_0[65]);
  nor NOR2_253 (KeyWire_0[136], N341, N659);
  xnor KeyGate_0_136(N731, keyIn_0_136, KeyWire_0[136]);
  nand NAND2_254 (KeyWire_0[137], N654, N261);
  xnor KeyGate_0_137(KeyNOTWire_0[66], keyIn_0_137, KeyWire_0[137]);
  not KeyNOTGate_0_66(N732, KeyNOTWire_0[66]);
  nand NAND3_255 (KeyWire_0[138], N644, N654, N261);
  xnor KeyGate_0_138(N733, keyIn_0_138, KeyWire_0[138]);
  nand NAND4_256 (KeyWire_0[139], N635, N644, N654, N261);
  xor KeyGate_0_139(KeyNOTWire_0[67], keyIn_0_139, KeyWire_0[139]);
  not KeyNOTGate_0_67(N734, KeyNOTWire_0[67]);
  not NOT1_257 (KeyWire_0[140], N662);
  xnor KeyGate_0_140(N735, keyIn_0_140, KeyWire_0[140]);
  and AND2_258 (KeyWire_0[141], N228, N665);
  xnor KeyGate_0_141(KeyNOTWire_0[68], keyIn_0_141, KeyWire_0[141]);
  not KeyNOTGate_0_68(N736, KeyNOTWire_0[68]);
  and AND2_259 (KeyWire_0[142], N237, N662);
  xor KeyGate_0_142(N737, keyIn_0_142, KeyWire_0[142]);
  not NOT1_260 (KeyWire_0[143], N670);
  xor KeyGate_0_143(N738, keyIn_0_143, KeyWire_0[143]);
  and AND2_261 (KeyWire_0[144], N228, N673);
  xor KeyGate_0_144(N739, keyIn_0_144, KeyWire_0[144]);
  and AND2_262 (KeyWire_0[145], N237, N670);
  xor KeyGate_0_145(N740, keyIn_0_145, KeyWire_0[145]);
  not NOT1_263 (KeyWire_0[146], N678);
  xor KeyGate_0_146(KeyNOTWire_0[69], keyIn_0_146, KeyWire_0[146]);
  not KeyNOTGate_0_69(N741, KeyNOTWire_0[69]);
  and AND2_264 (KeyWire_0[147], N228, N682);
  xnor KeyGate_0_147(KeyNOTWire_0[70], keyIn_0_147, KeyWire_0[147]);
  not KeyNOTGate_0_70(N742, KeyNOTWire_0[70]);
  and AND2_265 (KeyWire_0[148], N237, N678);
  xor KeyGate_0_148(N743, keyIn_0_148, KeyWire_0[148]);
  not NOT1_266 (KeyWire_0[149], N687);
  xnor KeyGate_0_149(KeyNOTWire_0[71], keyIn_0_149, KeyWire_0[149]);
  not KeyNOTGate_0_71(N744, KeyNOTWire_0[71]);
  and AND2_267 (KeyWire_0[150], N228, N692);
  xnor KeyGate_0_150(N745, keyIn_0_150, KeyWire_0[150]);
  and AND2_268 (KeyWire_0[151], N237, N687);
  xnor KeyGate_0_151(KeyNOTWire_0[72], keyIn_0_151, KeyWire_0[151]);
  not KeyNOTGate_0_72(N746, KeyNOTWire_0[72]);
  not NOT1_269 (KeyWire_0[152], N697);
  xor KeyGate_0_152(N747, keyIn_0_152, KeyWire_0[152]);
  and AND2_270 (KeyWire_0[153], N228, N700);
  xnor KeyGate_0_153(KeyNOTWire_0[73], keyIn_0_153, KeyWire_0[153]);
  not KeyNOTGate_0_73(N748, KeyNOTWire_0[73]);
  and AND2_271 (KeyWire_0[154], N237, N697);
  xor KeyGate_0_154(KeyNOTWire_0[74], keyIn_0_154, KeyWire_0[154]);
  not KeyNOTGate_0_74(N749, KeyNOTWire_0[74]);
  not NOT1_272 (KeyWire_0[155], N705);
  xnor KeyGate_0_155(KeyNOTWire_0[75], keyIn_0_155, KeyWire_0[155]);
  not KeyNOTGate_0_75(N750, KeyNOTWire_0[75]);
  and AND2_273 (KeyWire_0[156], N228, N708);
  xnor KeyGate_0_156(KeyNOTWire_0[76], keyIn_0_156, KeyWire_0[156]);
  not KeyNOTGate_0_76(N751, KeyNOTWire_0[76]);
  and AND2_274 (KeyWire_0[157], N237, N705);
  xnor KeyGate_0_157(KeyNOTWire_0[77], keyIn_0_157, KeyWire_0[157]);
  not KeyNOTGate_0_77(N752, KeyNOTWire_0[77]);
  not NOT1_275 (KeyWire_0[158], N713);
  xnor KeyGate_0_158(KeyNOTWire_0[78], keyIn_0_158, KeyWire_0[158]);
  not KeyNOTGate_0_78(N753, KeyNOTWire_0[78]);
  and AND2_276 (KeyWire_0[159], N228, N717);
  xnor KeyGate_0_159(KeyNOTWire_0[79], keyIn_0_159, KeyWire_0[159]);
  not KeyNOTGate_0_79(N754, KeyNOTWire_0[79]);
  and AND2_277 (KeyWire_0[160], N237, N713);
  xor KeyGate_0_160(KeyNOTWire_0[80], keyIn_0_160, KeyWire_0[160]);
  not KeyNOTGate_0_80(N755, KeyNOTWire_0[80]);
  not NOT1_278 (KeyWire_0[161], N722);
  xor KeyGate_0_161(KeyNOTWire_0[81], keyIn_0_161, KeyWire_0[161]);
  not KeyNOTGate_0_81(N756, KeyNOTWire_0[81]);
  nor NOR2_279 (KeyWire_0[162], N727, N261);
  xnor KeyGate_0_162(N757, keyIn_0_162, KeyWire_0[162]);
  and AND2_280 (KeyWire_0[163], N727, N261);
  xnor KeyGate_0_163(N758, keyIn_0_163, KeyWire_0[163]);
  and AND2_281 (KeyWire_0[164], N228, N727);
  xnor KeyGate_0_164(N759, keyIn_0_164, KeyWire_0[164]);
  and AND2_282 (KeyWire_0[165], N237, N722);
  xnor KeyGate_0_165(N760, keyIn_0_165, KeyWire_0[165]);
  nand NAND2_283 (KeyWire_0[166], N644, N722);
  xor KeyGate_0_166(N761, keyIn_0_166, KeyWire_0[166]);
  nand NAND2_284 (KeyWire_0[167], N635, N713);
  xor KeyGate_0_167(N762, keyIn_0_167, KeyWire_0[167]);
  nand NAND3_285 (KeyWire_0[168], N635, N644, N722);
  xnor KeyGate_0_168(N763, keyIn_0_168, KeyWire_0[168]);
  nand NAND2_286 (KeyWire_0[169], N609, N687);
  xor KeyGate_0_169(KeyNOTWire_0[82], keyIn_0_169, KeyWire_0[169]);
  not KeyNOTGate_0_82(N764, KeyNOTWire_0[82]);
  nand NAND2_287 (KeyWire_0[170], N600, N678);
  xor KeyGate_0_170(KeyNOTWire_0[83], keyIn_0_170, KeyWire_0[170]);
  not KeyNOTGate_0_83(N765, KeyNOTWire_0[83]);
  nand NAND3_288 (KeyWire_0[171], N600, N609, N687);
  xor KeyGate_0_171(KeyNOTWire_0[84], keyIn_0_171, KeyWire_0[171]);
  not KeyNOTGate_0_84(N766, KeyNOTWire_0[84]);
buf BUFF1_289 (N767, N660);
buf BUFF1_290 (N768, N661);
  nor NOR2_291 (KeyWire_0[172], N736, N737);
  xnor KeyGate_0_172(N769, keyIn_0_172, KeyWire_0[172]);
  nor NOR2_292 (KeyWire_0[173], N739, N740);
  xor KeyGate_0_173(KeyNOTWire_0[85], keyIn_0_173, KeyWire_0[173]);
  not KeyNOTGate_0_85(N770, KeyNOTWire_0[85]);
  nor NOR2_293 (KeyWire_0[174], N742, N743);
  xnor KeyGate_0_174(N771, keyIn_0_174, KeyWire_0[174]);
  nor NOR2_294 (KeyWire_0[175], N745, N746);
  xnor KeyGate_0_175(N772, keyIn_0_175, KeyWire_0[175]);
  nand NAND4_295 (KeyWire_0[176], N750, N762, N763, N734);
  xnor KeyGate_0_176(N773, keyIn_0_176, KeyWire_0[176]);
  nor NOR2_296 (KeyWire_0[177], N748, N749);
  xnor KeyGate_0_177(KeyNOTWire_0[86], keyIn_0_177, KeyWire_0[177]);
  not KeyNOTGate_0_86(N777, KeyNOTWire_0[86]);
  nand NAND3_297 (KeyWire_0[178], N753, N761, N733);
  xnor KeyGate_0_178(KeyNOTWire_0[87], keyIn_0_178, KeyWire_0[178]);
  not KeyNOTGate_0_87(N778, KeyNOTWire_0[87]);
  nor NOR2_298 (KeyWire_0[179], N751, N752);
  xnor KeyGate_0_179(N781, keyIn_0_179, KeyWire_0[179]);
  nand NAND2_299 (KeyWire_0[180], N756, N732);
  xor KeyGate_0_180(KeyNOTWire_0[88], keyIn_0_180, KeyWire_0[180]);
  not KeyNOTGate_0_88(N782, KeyNOTWire_0[88]);
  nor NOR2_300 (KeyWire_0[181], N754, N755);
  xor KeyGate_0_181(KeyNOTWire_0[89], keyIn_0_181, KeyWire_0[181]);
  not KeyNOTGate_0_89(N785, KeyNOTWire_0[89]);
  nor NOR2_301 (KeyWire_0[182], N757, N758);
  xnor KeyGate_0_182(N786, keyIn_0_182, KeyWire_0[182]);
  nor NOR2_302 (KeyWire_0[183], N759, N760);
  xnor KeyGate_0_183(N787, keyIn_0_183, KeyWire_0[183]);
  nor NOR2_303 (KeyWire_0[184], N700, N773);
  xnor KeyGate_0_184(KeyNOTWire_0[90], keyIn_0_184, KeyWire_0[184]);
  not KeyNOTGate_0_90(N788, KeyNOTWire_0[90]);
  and AND2_304 (KeyWire_0[185], N700, N773);
  xor KeyGate_0_185(KeyNOTWire_0[91], keyIn_0_185, KeyWire_0[185]);
  not KeyNOTGate_0_91(N789, KeyNOTWire_0[91]);
  nor NOR2_305 (KeyWire_0[186], N708, N778);
  xnor KeyGate_0_186(KeyNOTWire_0[92], keyIn_0_186, KeyWire_0[186]);
  not KeyNOTGate_0_92(N790, KeyNOTWire_0[92]);
  and AND2_306 (KeyWire_0[187], N708, N778);
  xor KeyGate_0_187(N791, keyIn_0_187, KeyWire_0[187]);
  nor NOR2_307 (KeyWire_0[188], N717, N782);
  xnor KeyGate_0_188(KeyNOTWire_0[93], keyIn_0_188, KeyWire_0[188]);
  not KeyNOTGate_0_93(N792, KeyNOTWire_0[93]);
  and AND2_308 (KeyWire_0[189], N717, N782);
  xor KeyGate_0_189(N793, keyIn_0_189, KeyWire_0[189]);
  and AND2_309 (KeyWire_0[190], N219, N786);
  xnor KeyGate_0_190(N794, keyIn_0_190, KeyWire_0[190]);
  nand NAND2_310 (KeyWire_0[191], N628, N773);
  xnor KeyGate_0_191(N795, keyIn_0_191, KeyWire_0[191]);
  nand NAND2_311 (KeyWire_0[192], N795, N747);
  xor KeyGate_0_192(N796, keyIn_0_192, KeyWire_0[192]);
  nor NOR2_312 (KeyWire_0[193], N788, N789);
  xnor KeyGate_0_193(N802, keyIn_0_193, KeyWire_0[193]);
  nor NOR2_313 (KeyWire_0[194], N790, N791);
  xnor KeyGate_0_194(N803, keyIn_0_194, KeyWire_0[194]);
  nor NOR2_314 (KeyWire_0[195], N792, N793);
  xnor KeyGate_0_195(N804, keyIn_0_195, KeyWire_0[195]);
  nor NOR2_315 (KeyWire_0[196], N340, N794);
  xnor KeyGate_0_196(N805, keyIn_0_196, KeyWire_0[196]);
  nor NOR2_316 (KeyWire_0[197], N692, N796);
  xor KeyGate_0_197(N806, keyIn_0_197, KeyWire_0[197]);
  and AND2_317 (KeyWire_0[198], N692, N796);
  xnor KeyGate_0_198(KeyNOTWire_0[94], keyIn_0_198, KeyWire_0[198]);
  not KeyNOTGate_0_94(N807, KeyNOTWire_0[94]);
  and AND2_318 (KeyWire_0[199], N219, N802);
  xnor KeyGate_0_199(KeyNOTWire_0[95], keyIn_0_199, KeyWire_0[199]);
  not KeyNOTGate_0_95(N808, KeyNOTWire_0[95]);
  and AND2_319 (KeyWire_0[200], N219, N803);
  xor KeyGate_0_200(KeyNOTWire_0[96], keyIn_0_200, KeyWire_0[200]);
  not KeyNOTGate_0_96(N809, KeyNOTWire_0[96]);
  and AND2_320 (KeyWire_0[201], N219, N804);
  xnor KeyGate_0_201(N810, keyIn_0_201, KeyWire_0[201]);
  nand NAND4_321 (KeyWire_0[202], N805, N787, N731, N529);
  xor KeyGate_0_202(N811, keyIn_0_202, KeyWire_0[202]);
  nand NAND2_322 (KeyWire_0[203], N619, N796);
  xnor KeyGate_0_203(KeyNOTWire_0[97], keyIn_0_203, KeyWire_0[203]);
  not KeyNOTGate_0_97(N812, KeyNOTWire_0[97]);
  nand NAND3_323 (KeyWire_0[204], N609, N619, N796);
  xnor KeyGate_0_204(KeyNOTWire_0[98], keyIn_0_204, KeyWire_0[204]);
  not KeyNOTGate_0_98(N813, KeyNOTWire_0[98]);
  nand NAND4_324 (KeyWire_0[205], N600, N609, N619, N796);
  xnor KeyGate_0_205(N814, keyIn_0_205, KeyWire_0[205]);
  nand NAND4_325 (KeyWire_0[206], N738, N765, N766, N814);
  xnor KeyGate_0_206(KeyNOTWire_0[99], keyIn_0_206, KeyWire_0[206]);
  not KeyNOTGate_0_99(N815, KeyNOTWire_0[99]);
  nand NAND3_326 (KeyWire_0[207], N741, N764, N813);
  xnor KeyGate_0_207(N819, keyIn_0_207, KeyWire_0[207]);
  nand NAND2_327 (KeyWire_0[208], N744, N812);
  xor KeyGate_0_208(N822, keyIn_0_208, KeyWire_0[208]);
  nor NOR2_328 (KeyWire_0[209], N806, N807);
  xnor KeyGate_0_209(KeyNOTWire_0[100], keyIn_0_209, KeyWire_0[209]);
  not KeyNOTGate_0_100(N825, KeyNOTWire_0[100]);
  nor NOR2_329 (KeyWire_0[210], N335, N808);
  xor KeyGate_0_210(N826, keyIn_0_210, KeyWire_0[210]);
  nor NOR2_330 (KeyWire_0[211], N336, N809);
  xor KeyGate_0_211(N827, keyIn_0_211, KeyWire_0[211]);
  nor NOR2_331 (KeyWire_0[212], N338, N810);
  xnor KeyGate_0_212(KeyNOTWire_0[101], keyIn_0_212, KeyWire_0[212]);
  not KeyNOTGate_0_101(N828, KeyNOTWire_0[101]);
  not NOT1_332 (KeyWire_0[213], N811);
  xnor KeyGate_0_213(KeyNOTWire_0[102], keyIn_0_213, KeyWire_0[213]);
  not KeyNOTGate_0_102(N829, KeyNOTWire_0[102]);
  nor NOR2_333 (KeyWire_0[214], N665, N815);
  xor KeyGate_0_214(N830, keyIn_0_214, KeyWire_0[214]);
  and AND2_334 (KeyWire_0[215], N665, N815);
  xor KeyGate_0_215(N831, keyIn_0_215, KeyWire_0[215]);
  nor NOR2_335 (KeyWire_0[216], N673, N819);
  xor KeyGate_0_216(KeyNOTWire_0[103], keyIn_0_216, KeyWire_0[216]);
  not KeyNOTGate_0_103(N832, KeyNOTWire_0[103]);
  and AND2_336 (KeyWire_0[217], N673, N819);
  xnor KeyGate_0_217(N833, keyIn_0_217, KeyWire_0[217]);
  nor NOR2_337 (KeyWire_0[218], N682, N822);
  xor KeyGate_0_218(N834, keyIn_0_218, KeyWire_0[218]);
  and AND2_338 (KeyWire_0[219], N682, N822);
  xor KeyGate_0_219(KeyNOTWire_0[104], keyIn_0_219, KeyWire_0[219]);
  not KeyNOTGate_0_104(N835, KeyNOTWire_0[104]);
  and AND2_339 (KeyWire_0[220], N219, N825);
  xnor KeyGate_0_220(KeyNOTWire_0[105], keyIn_0_220, KeyWire_0[220]);
  not KeyNOTGate_0_105(N836, KeyNOTWire_0[105]);
  nand NAND3_340 (KeyWire_0[221], N826, N777, N704);
  xor KeyGate_0_221(KeyNOTWire_0[106], keyIn_0_221, KeyWire_0[221]);
  not KeyNOTGate_0_106(N837, KeyNOTWire_0[106]);
  nand NAND4_341 (KeyWire_0[222], N827, N781, N712, N527);
  xnor KeyGate_0_222(KeyNOTWire_0[107], keyIn_0_222, KeyWire_0[222]);
  not KeyNOTGate_0_107(N838, KeyNOTWire_0[107]);
  nand NAND4_342 (KeyWire_0[223], N828, N785, N721, N528);
  xnor KeyGate_0_223(KeyNOTWire_0[108], keyIn_0_223, KeyWire_0[223]);
  not KeyNOTGate_0_108(N839, KeyNOTWire_0[108]);
  not NOT1_343 (KeyWire_0[224], N829);
  xnor KeyGate_0_224(KeyNOTWire_0[109], keyIn_0_224, KeyWire_0[224]);
  not KeyNOTGate_0_109(N840, KeyNOTWire_0[109]);
  nand NAND2_344 (KeyWire_0[225], N815, N593);
  xor KeyGate_0_225(KeyNOTWire_0[110], keyIn_0_225, KeyWire_0[225]);
  not KeyNOTGate_0_110(N841, KeyNOTWire_0[110]);
  nor NOR2_345 (KeyWire_0[226], N830, N831);
  xor KeyGate_0_226(KeyNOTWire_0[111], keyIn_0_226, KeyWire_0[226]);
  not KeyNOTGate_0_111(N842, KeyNOTWire_0[111]);
  nor NOR2_346 (KeyWire_0[227], N832, N833);
  xor KeyGate_0_227(N843, keyIn_0_227, KeyWire_0[227]);
  nor NOR2_347 (KeyWire_0[228], N834, N835);
  xnor KeyGate_0_228(KeyNOTWire_0[112], keyIn_0_228, KeyWire_0[228]);
  not KeyNOTGate_0_112(N844, KeyNOTWire_0[112]);
  nor NOR2_348 (KeyWire_0[229], N334, N836);
  xor KeyGate_0_229(KeyNOTWire_0[113], keyIn_0_229, KeyWire_0[229]);
  not KeyNOTGate_0_113(N845, KeyNOTWire_0[113]);
  not NOT1_349 (KeyWire_0[230], N837);
  xnor KeyGate_0_230(KeyNOTWire_0[114], keyIn_0_230, KeyWire_0[230]);
  not KeyNOTGate_0_114(N846, KeyNOTWire_0[114]);
  not NOT1_350 (KeyWire_0[231], N838);
  xnor KeyGate_0_231(N847, keyIn_0_231, KeyWire_0[231]);
  not NOT1_351 (KeyWire_0[232], N839);
  xnor KeyGate_0_232(KeyNOTWire_0[115], keyIn_0_232, KeyWire_0[232]);
  not KeyNOTGate_0_115(N848, KeyNOTWire_0[115]);
  and AND2_352 (KeyWire_0[233], N735, N841);
  xor KeyGate_0_233(KeyNOTWire_0[116], keyIn_0_233, KeyWire_0[233]);
  not KeyNOTGate_0_116(N849, KeyNOTWire_0[116]);
buf BUFF1_353 (N850, N840);
  and AND2_354 (KeyWire_0[234], N219, N842);
  xor KeyGate_0_234(N851, keyIn_0_234, KeyWire_0[234]);
  and AND2_355 (KeyWire_0[235], N219, N843);
  xnor KeyGate_0_235(N852, keyIn_0_235, KeyWire_0[235]);
  and AND2_356 (KeyWire_0[236], N219, N844);
  xor KeyGate_0_236(N853, keyIn_0_236, KeyWire_0[236]);
  nand NAND3_357 (KeyWire_0[237], N845, N772, N696);
  xnor KeyGate_0_237(N854, keyIn_0_237, KeyWire_0[237]);
  not NOT1_358 (KeyWire_0[238], N846);
  xor KeyGate_0_238(N855, keyIn_0_238, KeyWire_0[238]);
  not NOT1_359 (KeyWire_0[239], N847);
  xor KeyGate_0_239(KeyNOTWire_0[117], keyIn_0_239, KeyWire_0[239]);
  not KeyNOTGate_0_117(N856, KeyNOTWire_0[117]);
  not NOT1_360 (KeyWire_0[240], N848);
  xor KeyGate_0_240(N857, keyIn_0_240, KeyWire_0[240]);
  not NOT1_361 (KeyWire_0[241], N849);
  xor KeyGate_0_241(N858, keyIn_0_241, KeyWire_0[241]);
  nor NOR2_362 (KeyWire_0[242], N417, N851);
  xor KeyGate_0_242(N859, keyIn_0_242, KeyWire_0[242]);
  nor NOR2_363 (KeyWire_0[243], N332, N852);
  xnor KeyGate_0_243(KeyNOTWire_0[118], keyIn_0_243, KeyWire_0[243]);
  not KeyNOTGate_0_118(N860, KeyNOTWire_0[118]);
  nor NOR2_364 (KeyWire_0[244], N333, N853);
  xor KeyGate_0_244(KeyNOTWire_0[119], keyIn_0_244, KeyWire_0[244]);
  not KeyNOTGate_0_119(N861, KeyNOTWire_0[119]);
  not NOT1_365 (KeyWire_0[245], N854);
  xnor KeyGate_0_245(KeyNOTWire_0[120], keyIn_0_245, KeyWire_0[245]);
  not KeyNOTGate_0_120(N862, KeyNOTWire_0[120]);
buf BUFF1_366 (N863, N855);
buf BUFF1_367 (N864, N856);
buf BUFF1_368 (N865, N857);
buf BUFF1_369 (N866, N858);
  nand NAND3_370 (KeyWire_0[246], N859, N769, N669);
  xnor KeyGate_0_246(N867, keyIn_0_246, KeyWire_0[246]);
  nand NAND3_371 (KeyWire_0[247], N860, N770, N677);
  xnor KeyGate_0_247(N868, keyIn_0_247, KeyWire_0[247]);
  nand NAND3_372 (KeyWire_0[248], N861, N771, N686);
  xor KeyGate_0_248(KeyNOTWire_0[121], keyIn_0_248, KeyWire_0[248]);
  not KeyNOTGate_0_121(N869, KeyNOTWire_0[121]);
  not NOT1_373 (KeyWire_0[249], N862);
  xor KeyGate_0_249(KeyNOTWire_0[122], keyIn_0_249, KeyWire_0[249]);
  not KeyNOTGate_0_122(N870, KeyNOTWire_0[122]);
  not NOT1_374 (KeyWire_0[250], N867);
  xnor KeyGate_0_250(N871, keyIn_0_250, KeyWire_0[250]);
  not NOT1_375 (KeyWire_0[251], N868);
  xnor KeyGate_0_251(KeyNOTWire_0[123], keyIn_0_251, KeyWire_0[251]);
  not KeyNOTGate_0_123(N872, KeyNOTWire_0[123]);
  not NOT1_376 (KeyWire_0[252], N869);
  xor KeyGate_0_252(N873, keyIn_0_252, KeyWire_0[252]);
buf BUFF1_377 (N874, N870);
  not NOT1_378 (KeyWire_0[253], N871);
  xor KeyGate_0_253(N875, keyIn_0_253, KeyWire_0[253]);
  not NOT1_379 (KeyWire_0[254], N872);
  xnor KeyGate_0_254(KeyNOTWire_0[124], keyIn_0_254, KeyWire_0[254]);
  not KeyNOTGate_0_124(N876, KeyNOTWire_0[124]);
  not NOT1_380 (KeyWire_0[255], N873);
  xor KeyGate_0_255(KeyNOTWire_0[125], keyIn_0_255, KeyWire_0[255]);
  not KeyNOTGate_0_125(N877, KeyNOTWire_0[125]);
buf BUFF1_381 (N878, N875);
buf BUFF1_382 (N879, N876);
buf BUFF1_383 (N880, N877);

endmodule
